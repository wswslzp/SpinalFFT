// Generator : SpinalHDL v1.4.1    git head : 99d6d471af204b6d7d9f63fae58757e9d3c7b944
// Component : MyFFT



module MyFFT (
  input               io_data_in_valid,
  input      [15:0]   io_data_in_payload_0_real,
  input      [15:0]   io_data_in_payload_0_imag,
  input      [15:0]   io_data_in_payload_1_real,
  input      [15:0]   io_data_in_payload_1_imag,
  input      [15:0]   io_data_in_payload_2_real,
  input      [15:0]   io_data_in_payload_2_imag,
  input      [15:0]   io_data_in_payload_3_real,
  input      [15:0]   io_data_in_payload_3_imag,
  input      [15:0]   io_data_in_payload_4_real,
  input      [15:0]   io_data_in_payload_4_imag,
  input      [15:0]   io_data_in_payload_5_real,
  input      [15:0]   io_data_in_payload_5_imag,
  input      [15:0]   io_data_in_payload_6_real,
  input      [15:0]   io_data_in_payload_6_imag,
  input      [15:0]   io_data_in_payload_7_real,
  input      [15:0]   io_data_in_payload_7_imag,
  input      [15:0]   io_data_in_payload_8_real,
  input      [15:0]   io_data_in_payload_8_imag,
  input      [15:0]   io_data_in_payload_9_real,
  input      [15:0]   io_data_in_payload_9_imag,
  input      [15:0]   io_data_in_payload_10_real,
  input      [15:0]   io_data_in_payload_10_imag,
  input      [15:0]   io_data_in_payload_11_real,
  input      [15:0]   io_data_in_payload_11_imag,
  input      [15:0]   io_data_in_payload_12_real,
  input      [15:0]   io_data_in_payload_12_imag,
  input      [15:0]   io_data_in_payload_13_real,
  input      [15:0]   io_data_in_payload_13_imag,
  input      [15:0]   io_data_in_payload_14_real,
  input      [15:0]   io_data_in_payload_14_imag,
  input      [15:0]   io_data_in_payload_15_real,
  input      [15:0]   io_data_in_payload_15_imag,
  input      [15:0]   io_data_in_payload_16_real,
  input      [15:0]   io_data_in_payload_16_imag,
  input      [15:0]   io_data_in_payload_17_real,
  input      [15:0]   io_data_in_payload_17_imag,
  input      [15:0]   io_data_in_payload_18_real,
  input      [15:0]   io_data_in_payload_18_imag,
  input      [15:0]   io_data_in_payload_19_real,
  input      [15:0]   io_data_in_payload_19_imag,
  input      [15:0]   io_data_in_payload_20_real,
  input      [15:0]   io_data_in_payload_20_imag,
  input      [15:0]   io_data_in_payload_21_real,
  input      [15:0]   io_data_in_payload_21_imag,
  input      [15:0]   io_data_in_payload_22_real,
  input      [15:0]   io_data_in_payload_22_imag,
  input      [15:0]   io_data_in_payload_23_real,
  input      [15:0]   io_data_in_payload_23_imag,
  input      [15:0]   io_data_in_payload_24_real,
  input      [15:0]   io_data_in_payload_24_imag,
  input      [15:0]   io_data_in_payload_25_real,
  input      [15:0]   io_data_in_payload_25_imag,
  input      [15:0]   io_data_in_payload_26_real,
  input      [15:0]   io_data_in_payload_26_imag,
  input      [15:0]   io_data_in_payload_27_real,
  input      [15:0]   io_data_in_payload_27_imag,
  input      [15:0]   io_data_in_payload_28_real,
  input      [15:0]   io_data_in_payload_28_imag,
  input      [15:0]   io_data_in_payload_29_real,
  input      [15:0]   io_data_in_payload_29_imag,
  input      [15:0]   io_data_in_payload_30_real,
  input      [15:0]   io_data_in_payload_30_imag,
  input      [15:0]   io_data_in_payload_31_real,
  input      [15:0]   io_data_in_payload_31_imag,
  input      [15:0]   io_data_in_payload_32_real,
  input      [15:0]   io_data_in_payload_32_imag,
  input      [15:0]   io_data_in_payload_33_real,
  input      [15:0]   io_data_in_payload_33_imag,
  input      [15:0]   io_data_in_payload_34_real,
  input      [15:0]   io_data_in_payload_34_imag,
  input      [15:0]   io_data_in_payload_35_real,
  input      [15:0]   io_data_in_payload_35_imag,
  input      [15:0]   io_data_in_payload_36_real,
  input      [15:0]   io_data_in_payload_36_imag,
  input      [15:0]   io_data_in_payload_37_real,
  input      [15:0]   io_data_in_payload_37_imag,
  input      [15:0]   io_data_in_payload_38_real,
  input      [15:0]   io_data_in_payload_38_imag,
  input      [15:0]   io_data_in_payload_39_real,
  input      [15:0]   io_data_in_payload_39_imag,
  input      [15:0]   io_data_in_payload_40_real,
  input      [15:0]   io_data_in_payload_40_imag,
  input      [15:0]   io_data_in_payload_41_real,
  input      [15:0]   io_data_in_payload_41_imag,
  input      [15:0]   io_data_in_payload_42_real,
  input      [15:0]   io_data_in_payload_42_imag,
  input      [15:0]   io_data_in_payload_43_real,
  input      [15:0]   io_data_in_payload_43_imag,
  input      [15:0]   io_data_in_payload_44_real,
  input      [15:0]   io_data_in_payload_44_imag,
  input      [15:0]   io_data_in_payload_45_real,
  input      [15:0]   io_data_in_payload_45_imag,
  input      [15:0]   io_data_in_payload_46_real,
  input      [15:0]   io_data_in_payload_46_imag,
  input      [15:0]   io_data_in_payload_47_real,
  input      [15:0]   io_data_in_payload_47_imag,
  input      [15:0]   io_data_in_payload_48_real,
  input      [15:0]   io_data_in_payload_48_imag,
  input      [15:0]   io_data_in_payload_49_real,
  input      [15:0]   io_data_in_payload_49_imag,
  input      [15:0]   io_data_in_payload_50_real,
  input      [15:0]   io_data_in_payload_50_imag,
  input      [15:0]   io_data_in_payload_51_real,
  input      [15:0]   io_data_in_payload_51_imag,
  input      [15:0]   io_data_in_payload_52_real,
  input      [15:0]   io_data_in_payload_52_imag,
  input      [15:0]   io_data_in_payload_53_real,
  input      [15:0]   io_data_in_payload_53_imag,
  input      [15:0]   io_data_in_payload_54_real,
  input      [15:0]   io_data_in_payload_54_imag,
  input      [15:0]   io_data_in_payload_55_real,
  input      [15:0]   io_data_in_payload_55_imag,
  input      [15:0]   io_data_in_payload_56_real,
  input      [15:0]   io_data_in_payload_56_imag,
  input      [15:0]   io_data_in_payload_57_real,
  input      [15:0]   io_data_in_payload_57_imag,
  input      [15:0]   io_data_in_payload_58_real,
  input      [15:0]   io_data_in_payload_58_imag,
  input      [15:0]   io_data_in_payload_59_real,
  input      [15:0]   io_data_in_payload_59_imag,
  input      [15:0]   io_data_in_payload_60_real,
  input      [15:0]   io_data_in_payload_60_imag,
  input      [15:0]   io_data_in_payload_61_real,
  input      [15:0]   io_data_in_payload_61_imag,
  input      [15:0]   io_data_in_payload_62_real,
  input      [15:0]   io_data_in_payload_62_imag,
  input      [15:0]   io_data_in_payload_63_real,
  input      [15:0]   io_data_in_payload_63_imag,
  input      [15:0]   io_data_in_payload_64_real,
  input      [15:0]   io_data_in_payload_64_imag,
  input      [15:0]   io_data_in_payload_65_real,
  input      [15:0]   io_data_in_payload_65_imag,
  input      [15:0]   io_data_in_payload_66_real,
  input      [15:0]   io_data_in_payload_66_imag,
  input      [15:0]   io_data_in_payload_67_real,
  input      [15:0]   io_data_in_payload_67_imag,
  input      [15:0]   io_data_in_payload_68_real,
  input      [15:0]   io_data_in_payload_68_imag,
  input      [15:0]   io_data_in_payload_69_real,
  input      [15:0]   io_data_in_payload_69_imag,
  input      [15:0]   io_data_in_payload_70_real,
  input      [15:0]   io_data_in_payload_70_imag,
  input      [15:0]   io_data_in_payload_71_real,
  input      [15:0]   io_data_in_payload_71_imag,
  input      [15:0]   io_data_in_payload_72_real,
  input      [15:0]   io_data_in_payload_72_imag,
  input      [15:0]   io_data_in_payload_73_real,
  input      [15:0]   io_data_in_payload_73_imag,
  input      [15:0]   io_data_in_payload_74_real,
  input      [15:0]   io_data_in_payload_74_imag,
  input      [15:0]   io_data_in_payload_75_real,
  input      [15:0]   io_data_in_payload_75_imag,
  input      [15:0]   io_data_in_payload_76_real,
  input      [15:0]   io_data_in_payload_76_imag,
  input      [15:0]   io_data_in_payload_77_real,
  input      [15:0]   io_data_in_payload_77_imag,
  input      [15:0]   io_data_in_payload_78_real,
  input      [15:0]   io_data_in_payload_78_imag,
  input      [15:0]   io_data_in_payload_79_real,
  input      [15:0]   io_data_in_payload_79_imag,
  input      [15:0]   io_data_in_payload_80_real,
  input      [15:0]   io_data_in_payload_80_imag,
  input      [15:0]   io_data_in_payload_81_real,
  input      [15:0]   io_data_in_payload_81_imag,
  input      [15:0]   io_data_in_payload_82_real,
  input      [15:0]   io_data_in_payload_82_imag,
  input      [15:0]   io_data_in_payload_83_real,
  input      [15:0]   io_data_in_payload_83_imag,
  input      [15:0]   io_data_in_payload_84_real,
  input      [15:0]   io_data_in_payload_84_imag,
  input      [15:0]   io_data_in_payload_85_real,
  input      [15:0]   io_data_in_payload_85_imag,
  input      [15:0]   io_data_in_payload_86_real,
  input      [15:0]   io_data_in_payload_86_imag,
  input      [15:0]   io_data_in_payload_87_real,
  input      [15:0]   io_data_in_payload_87_imag,
  input      [15:0]   io_data_in_payload_88_real,
  input      [15:0]   io_data_in_payload_88_imag,
  input      [15:0]   io_data_in_payload_89_real,
  input      [15:0]   io_data_in_payload_89_imag,
  input      [15:0]   io_data_in_payload_90_real,
  input      [15:0]   io_data_in_payload_90_imag,
  input      [15:0]   io_data_in_payload_91_real,
  input      [15:0]   io_data_in_payload_91_imag,
  input      [15:0]   io_data_in_payload_92_real,
  input      [15:0]   io_data_in_payload_92_imag,
  input      [15:0]   io_data_in_payload_93_real,
  input      [15:0]   io_data_in_payload_93_imag,
  input      [15:0]   io_data_in_payload_94_real,
  input      [15:0]   io_data_in_payload_94_imag,
  input      [15:0]   io_data_in_payload_95_real,
  input      [15:0]   io_data_in_payload_95_imag,
  input      [15:0]   io_data_in_payload_96_real,
  input      [15:0]   io_data_in_payload_96_imag,
  input      [15:0]   io_data_in_payload_97_real,
  input      [15:0]   io_data_in_payload_97_imag,
  input      [15:0]   io_data_in_payload_98_real,
  input      [15:0]   io_data_in_payload_98_imag,
  input      [15:0]   io_data_in_payload_99_real,
  input      [15:0]   io_data_in_payload_99_imag,
  input      [15:0]   io_data_in_payload_100_real,
  input      [15:0]   io_data_in_payload_100_imag,
  input      [15:0]   io_data_in_payload_101_real,
  input      [15:0]   io_data_in_payload_101_imag,
  input      [15:0]   io_data_in_payload_102_real,
  input      [15:0]   io_data_in_payload_102_imag,
  input      [15:0]   io_data_in_payload_103_real,
  input      [15:0]   io_data_in_payload_103_imag,
  input      [15:0]   io_data_in_payload_104_real,
  input      [15:0]   io_data_in_payload_104_imag,
  input      [15:0]   io_data_in_payload_105_real,
  input      [15:0]   io_data_in_payload_105_imag,
  input      [15:0]   io_data_in_payload_106_real,
  input      [15:0]   io_data_in_payload_106_imag,
  input      [15:0]   io_data_in_payload_107_real,
  input      [15:0]   io_data_in_payload_107_imag,
  input      [15:0]   io_data_in_payload_108_real,
  input      [15:0]   io_data_in_payload_108_imag,
  input      [15:0]   io_data_in_payload_109_real,
  input      [15:0]   io_data_in_payload_109_imag,
  input      [15:0]   io_data_in_payload_110_real,
  input      [15:0]   io_data_in_payload_110_imag,
  input      [15:0]   io_data_in_payload_111_real,
  input      [15:0]   io_data_in_payload_111_imag,
  input      [15:0]   io_data_in_payload_112_real,
  input      [15:0]   io_data_in_payload_112_imag,
  input      [15:0]   io_data_in_payload_113_real,
  input      [15:0]   io_data_in_payload_113_imag,
  input      [15:0]   io_data_in_payload_114_real,
  input      [15:0]   io_data_in_payload_114_imag,
  input      [15:0]   io_data_in_payload_115_real,
  input      [15:0]   io_data_in_payload_115_imag,
  input      [15:0]   io_data_in_payload_116_real,
  input      [15:0]   io_data_in_payload_116_imag,
  input      [15:0]   io_data_in_payload_117_real,
  input      [15:0]   io_data_in_payload_117_imag,
  input      [15:0]   io_data_in_payload_118_real,
  input      [15:0]   io_data_in_payload_118_imag,
  input      [15:0]   io_data_in_payload_119_real,
  input      [15:0]   io_data_in_payload_119_imag,
  input      [15:0]   io_data_in_payload_120_real,
  input      [15:0]   io_data_in_payload_120_imag,
  input      [15:0]   io_data_in_payload_121_real,
  input      [15:0]   io_data_in_payload_121_imag,
  input      [15:0]   io_data_in_payload_122_real,
  input      [15:0]   io_data_in_payload_122_imag,
  input      [15:0]   io_data_in_payload_123_real,
  input      [15:0]   io_data_in_payload_123_imag,
  input      [15:0]   io_data_in_payload_124_real,
  input      [15:0]   io_data_in_payload_124_imag,
  input      [15:0]   io_data_in_payload_125_real,
  input      [15:0]   io_data_in_payload_125_imag,
  input      [15:0]   io_data_in_payload_126_real,
  input      [15:0]   io_data_in_payload_126_imag,
  input      [15:0]   io_data_in_payload_127_real,
  input      [15:0]   io_data_in_payload_127_imag,
  output              io_data_out_valid,
  output     [15:0]   io_data_out_payload_0_real,
  output     [15:0]   io_data_out_payload_0_imag,
  output     [15:0]   io_data_out_payload_1_real,
  output     [15:0]   io_data_out_payload_1_imag,
  output     [15:0]   io_data_out_payload_2_real,
  output     [15:0]   io_data_out_payload_2_imag,
  output     [15:0]   io_data_out_payload_3_real,
  output     [15:0]   io_data_out_payload_3_imag,
  output     [15:0]   io_data_out_payload_4_real,
  output     [15:0]   io_data_out_payload_4_imag,
  output     [15:0]   io_data_out_payload_5_real,
  output     [15:0]   io_data_out_payload_5_imag,
  output     [15:0]   io_data_out_payload_6_real,
  output     [15:0]   io_data_out_payload_6_imag,
  output     [15:0]   io_data_out_payload_7_real,
  output     [15:0]   io_data_out_payload_7_imag,
  output     [15:0]   io_data_out_payload_8_real,
  output     [15:0]   io_data_out_payload_8_imag,
  output     [15:0]   io_data_out_payload_9_real,
  output     [15:0]   io_data_out_payload_9_imag,
  output     [15:0]   io_data_out_payload_10_real,
  output     [15:0]   io_data_out_payload_10_imag,
  output     [15:0]   io_data_out_payload_11_real,
  output     [15:0]   io_data_out_payload_11_imag,
  output     [15:0]   io_data_out_payload_12_real,
  output     [15:0]   io_data_out_payload_12_imag,
  output     [15:0]   io_data_out_payload_13_real,
  output     [15:0]   io_data_out_payload_13_imag,
  output     [15:0]   io_data_out_payload_14_real,
  output     [15:0]   io_data_out_payload_14_imag,
  output     [15:0]   io_data_out_payload_15_real,
  output     [15:0]   io_data_out_payload_15_imag,
  output     [15:0]   io_data_out_payload_16_real,
  output     [15:0]   io_data_out_payload_16_imag,
  output     [15:0]   io_data_out_payload_17_real,
  output     [15:0]   io_data_out_payload_17_imag,
  output     [15:0]   io_data_out_payload_18_real,
  output     [15:0]   io_data_out_payload_18_imag,
  output     [15:0]   io_data_out_payload_19_real,
  output     [15:0]   io_data_out_payload_19_imag,
  output     [15:0]   io_data_out_payload_20_real,
  output     [15:0]   io_data_out_payload_20_imag,
  output     [15:0]   io_data_out_payload_21_real,
  output     [15:0]   io_data_out_payload_21_imag,
  output     [15:0]   io_data_out_payload_22_real,
  output     [15:0]   io_data_out_payload_22_imag,
  output     [15:0]   io_data_out_payload_23_real,
  output     [15:0]   io_data_out_payload_23_imag,
  output     [15:0]   io_data_out_payload_24_real,
  output     [15:0]   io_data_out_payload_24_imag,
  output     [15:0]   io_data_out_payload_25_real,
  output     [15:0]   io_data_out_payload_25_imag,
  output     [15:0]   io_data_out_payload_26_real,
  output     [15:0]   io_data_out_payload_26_imag,
  output     [15:0]   io_data_out_payload_27_real,
  output     [15:0]   io_data_out_payload_27_imag,
  output     [15:0]   io_data_out_payload_28_real,
  output     [15:0]   io_data_out_payload_28_imag,
  output     [15:0]   io_data_out_payload_29_real,
  output     [15:0]   io_data_out_payload_29_imag,
  output     [15:0]   io_data_out_payload_30_real,
  output     [15:0]   io_data_out_payload_30_imag,
  output     [15:0]   io_data_out_payload_31_real,
  output     [15:0]   io_data_out_payload_31_imag,
  output     [15:0]   io_data_out_payload_32_real,
  output     [15:0]   io_data_out_payload_32_imag,
  output     [15:0]   io_data_out_payload_33_real,
  output     [15:0]   io_data_out_payload_33_imag,
  output     [15:0]   io_data_out_payload_34_real,
  output     [15:0]   io_data_out_payload_34_imag,
  output     [15:0]   io_data_out_payload_35_real,
  output     [15:0]   io_data_out_payload_35_imag,
  output     [15:0]   io_data_out_payload_36_real,
  output     [15:0]   io_data_out_payload_36_imag,
  output     [15:0]   io_data_out_payload_37_real,
  output     [15:0]   io_data_out_payload_37_imag,
  output     [15:0]   io_data_out_payload_38_real,
  output     [15:0]   io_data_out_payload_38_imag,
  output     [15:0]   io_data_out_payload_39_real,
  output     [15:0]   io_data_out_payload_39_imag,
  output     [15:0]   io_data_out_payload_40_real,
  output     [15:0]   io_data_out_payload_40_imag,
  output     [15:0]   io_data_out_payload_41_real,
  output     [15:0]   io_data_out_payload_41_imag,
  output     [15:0]   io_data_out_payload_42_real,
  output     [15:0]   io_data_out_payload_42_imag,
  output     [15:0]   io_data_out_payload_43_real,
  output     [15:0]   io_data_out_payload_43_imag,
  output     [15:0]   io_data_out_payload_44_real,
  output     [15:0]   io_data_out_payload_44_imag,
  output     [15:0]   io_data_out_payload_45_real,
  output     [15:0]   io_data_out_payload_45_imag,
  output     [15:0]   io_data_out_payload_46_real,
  output     [15:0]   io_data_out_payload_46_imag,
  output     [15:0]   io_data_out_payload_47_real,
  output     [15:0]   io_data_out_payload_47_imag,
  output     [15:0]   io_data_out_payload_48_real,
  output     [15:0]   io_data_out_payload_48_imag,
  output     [15:0]   io_data_out_payload_49_real,
  output     [15:0]   io_data_out_payload_49_imag,
  output     [15:0]   io_data_out_payload_50_real,
  output     [15:0]   io_data_out_payload_50_imag,
  output     [15:0]   io_data_out_payload_51_real,
  output     [15:0]   io_data_out_payload_51_imag,
  output     [15:0]   io_data_out_payload_52_real,
  output     [15:0]   io_data_out_payload_52_imag,
  output     [15:0]   io_data_out_payload_53_real,
  output     [15:0]   io_data_out_payload_53_imag,
  output     [15:0]   io_data_out_payload_54_real,
  output     [15:0]   io_data_out_payload_54_imag,
  output     [15:0]   io_data_out_payload_55_real,
  output     [15:0]   io_data_out_payload_55_imag,
  output     [15:0]   io_data_out_payload_56_real,
  output     [15:0]   io_data_out_payload_56_imag,
  output     [15:0]   io_data_out_payload_57_real,
  output     [15:0]   io_data_out_payload_57_imag,
  output     [15:0]   io_data_out_payload_58_real,
  output     [15:0]   io_data_out_payload_58_imag,
  output     [15:0]   io_data_out_payload_59_real,
  output     [15:0]   io_data_out_payload_59_imag,
  output     [15:0]   io_data_out_payload_60_real,
  output     [15:0]   io_data_out_payload_60_imag,
  output     [15:0]   io_data_out_payload_61_real,
  output     [15:0]   io_data_out_payload_61_imag,
  output     [15:0]   io_data_out_payload_62_real,
  output     [15:0]   io_data_out_payload_62_imag,
  output     [15:0]   io_data_out_payload_63_real,
  output     [15:0]   io_data_out_payload_63_imag,
  output     [15:0]   io_data_out_payload_64_real,
  output     [15:0]   io_data_out_payload_64_imag,
  output     [15:0]   io_data_out_payload_65_real,
  output     [15:0]   io_data_out_payload_65_imag,
  output     [15:0]   io_data_out_payload_66_real,
  output     [15:0]   io_data_out_payload_66_imag,
  output     [15:0]   io_data_out_payload_67_real,
  output     [15:0]   io_data_out_payload_67_imag,
  output     [15:0]   io_data_out_payload_68_real,
  output     [15:0]   io_data_out_payload_68_imag,
  output     [15:0]   io_data_out_payload_69_real,
  output     [15:0]   io_data_out_payload_69_imag,
  output     [15:0]   io_data_out_payload_70_real,
  output     [15:0]   io_data_out_payload_70_imag,
  output     [15:0]   io_data_out_payload_71_real,
  output     [15:0]   io_data_out_payload_71_imag,
  output     [15:0]   io_data_out_payload_72_real,
  output     [15:0]   io_data_out_payload_72_imag,
  output     [15:0]   io_data_out_payload_73_real,
  output     [15:0]   io_data_out_payload_73_imag,
  output     [15:0]   io_data_out_payload_74_real,
  output     [15:0]   io_data_out_payload_74_imag,
  output     [15:0]   io_data_out_payload_75_real,
  output     [15:0]   io_data_out_payload_75_imag,
  output     [15:0]   io_data_out_payload_76_real,
  output     [15:0]   io_data_out_payload_76_imag,
  output     [15:0]   io_data_out_payload_77_real,
  output     [15:0]   io_data_out_payload_77_imag,
  output     [15:0]   io_data_out_payload_78_real,
  output     [15:0]   io_data_out_payload_78_imag,
  output     [15:0]   io_data_out_payload_79_real,
  output     [15:0]   io_data_out_payload_79_imag,
  output     [15:0]   io_data_out_payload_80_real,
  output     [15:0]   io_data_out_payload_80_imag,
  output     [15:0]   io_data_out_payload_81_real,
  output     [15:0]   io_data_out_payload_81_imag,
  output     [15:0]   io_data_out_payload_82_real,
  output     [15:0]   io_data_out_payload_82_imag,
  output     [15:0]   io_data_out_payload_83_real,
  output     [15:0]   io_data_out_payload_83_imag,
  output     [15:0]   io_data_out_payload_84_real,
  output     [15:0]   io_data_out_payload_84_imag,
  output     [15:0]   io_data_out_payload_85_real,
  output     [15:0]   io_data_out_payload_85_imag,
  output     [15:0]   io_data_out_payload_86_real,
  output     [15:0]   io_data_out_payload_86_imag,
  output     [15:0]   io_data_out_payload_87_real,
  output     [15:0]   io_data_out_payload_87_imag,
  output     [15:0]   io_data_out_payload_88_real,
  output     [15:0]   io_data_out_payload_88_imag,
  output     [15:0]   io_data_out_payload_89_real,
  output     [15:0]   io_data_out_payload_89_imag,
  output     [15:0]   io_data_out_payload_90_real,
  output     [15:0]   io_data_out_payload_90_imag,
  output     [15:0]   io_data_out_payload_91_real,
  output     [15:0]   io_data_out_payload_91_imag,
  output     [15:0]   io_data_out_payload_92_real,
  output     [15:0]   io_data_out_payload_92_imag,
  output     [15:0]   io_data_out_payload_93_real,
  output     [15:0]   io_data_out_payload_93_imag,
  output     [15:0]   io_data_out_payload_94_real,
  output     [15:0]   io_data_out_payload_94_imag,
  output     [15:0]   io_data_out_payload_95_real,
  output     [15:0]   io_data_out_payload_95_imag,
  output     [15:0]   io_data_out_payload_96_real,
  output     [15:0]   io_data_out_payload_96_imag,
  output     [15:0]   io_data_out_payload_97_real,
  output     [15:0]   io_data_out_payload_97_imag,
  output     [15:0]   io_data_out_payload_98_real,
  output     [15:0]   io_data_out_payload_98_imag,
  output     [15:0]   io_data_out_payload_99_real,
  output     [15:0]   io_data_out_payload_99_imag,
  output     [15:0]   io_data_out_payload_100_real,
  output     [15:0]   io_data_out_payload_100_imag,
  output     [15:0]   io_data_out_payload_101_real,
  output     [15:0]   io_data_out_payload_101_imag,
  output     [15:0]   io_data_out_payload_102_real,
  output     [15:0]   io_data_out_payload_102_imag,
  output     [15:0]   io_data_out_payload_103_real,
  output     [15:0]   io_data_out_payload_103_imag,
  output     [15:0]   io_data_out_payload_104_real,
  output     [15:0]   io_data_out_payload_104_imag,
  output     [15:0]   io_data_out_payload_105_real,
  output     [15:0]   io_data_out_payload_105_imag,
  output     [15:0]   io_data_out_payload_106_real,
  output     [15:0]   io_data_out_payload_106_imag,
  output     [15:0]   io_data_out_payload_107_real,
  output     [15:0]   io_data_out_payload_107_imag,
  output     [15:0]   io_data_out_payload_108_real,
  output     [15:0]   io_data_out_payload_108_imag,
  output     [15:0]   io_data_out_payload_109_real,
  output     [15:0]   io_data_out_payload_109_imag,
  output     [15:0]   io_data_out_payload_110_real,
  output     [15:0]   io_data_out_payload_110_imag,
  output     [15:0]   io_data_out_payload_111_real,
  output     [15:0]   io_data_out_payload_111_imag,
  output     [15:0]   io_data_out_payload_112_real,
  output     [15:0]   io_data_out_payload_112_imag,
  output     [15:0]   io_data_out_payload_113_real,
  output     [15:0]   io_data_out_payload_113_imag,
  output     [15:0]   io_data_out_payload_114_real,
  output     [15:0]   io_data_out_payload_114_imag,
  output     [15:0]   io_data_out_payload_115_real,
  output     [15:0]   io_data_out_payload_115_imag,
  output     [15:0]   io_data_out_payload_116_real,
  output     [15:0]   io_data_out_payload_116_imag,
  output     [15:0]   io_data_out_payload_117_real,
  output     [15:0]   io_data_out_payload_117_imag,
  output     [15:0]   io_data_out_payload_118_real,
  output     [15:0]   io_data_out_payload_118_imag,
  output     [15:0]   io_data_out_payload_119_real,
  output     [15:0]   io_data_out_payload_119_imag,
  output     [15:0]   io_data_out_payload_120_real,
  output     [15:0]   io_data_out_payload_120_imag,
  output     [15:0]   io_data_out_payload_121_real,
  output     [15:0]   io_data_out_payload_121_imag,
  output     [15:0]   io_data_out_payload_122_real,
  output     [15:0]   io_data_out_payload_122_imag,
  output     [15:0]   io_data_out_payload_123_real,
  output     [15:0]   io_data_out_payload_123_imag,
  output     [15:0]   io_data_out_payload_124_real,
  output     [15:0]   io_data_out_payload_124_imag,
  output     [15:0]   io_data_out_payload_125_real,
  output     [15:0]   io_data_out_payload_125_imag,
  output     [15:0]   io_data_out_payload_126_real,
  output     [15:0]   io_data_out_payload_126_imag,
  output     [15:0]   io_data_out_payload_127_real,
  output     [15:0]   io_data_out_payload_127_imag,
  input               clk,
  input               reset
);
  wire       [31:0]   _zz_1793;
  wire       [31:0]   _zz_1794;
  wire       [31:0]   _zz_1795;
  wire       [31:0]   _zz_1796;
  wire       [31:0]   _zz_1797;
  wire       [31:0]   _zz_1798;
  wire       [31:0]   _zz_1799;
  wire       [31:0]   _zz_1800;
  wire       [31:0]   _zz_1801;
  wire       [31:0]   _zz_1802;
  wire       [31:0]   _zz_1803;
  wire       [31:0]   _zz_1804;
  wire       [31:0]   _zz_1805;
  wire       [31:0]   _zz_1806;
  wire       [31:0]   _zz_1807;
  wire       [31:0]   _zz_1808;
  wire       [31:0]   _zz_1809;
  wire       [31:0]   _zz_1810;
  wire       [31:0]   _zz_1811;
  wire       [31:0]   _zz_1812;
  wire       [31:0]   _zz_1813;
  wire       [31:0]   _zz_1814;
  wire       [31:0]   _zz_1815;
  wire       [31:0]   _zz_1816;
  wire       [31:0]   _zz_1817;
  wire       [31:0]   _zz_1818;
  wire       [31:0]   _zz_1819;
  wire       [31:0]   _zz_1820;
  wire       [31:0]   _zz_1821;
  wire       [31:0]   _zz_1822;
  wire       [31:0]   _zz_1823;
  wire       [31:0]   _zz_1824;
  wire       [31:0]   _zz_1825;
  wire       [31:0]   _zz_1826;
  wire       [31:0]   _zz_1827;
  wire       [31:0]   _zz_1828;
  wire       [31:0]   _zz_1829;
  wire       [31:0]   _zz_1830;
  wire       [31:0]   _zz_1831;
  wire       [31:0]   _zz_1832;
  wire       [31:0]   _zz_1833;
  wire       [31:0]   _zz_1834;
  wire       [31:0]   _zz_1835;
  wire       [31:0]   _zz_1836;
  wire       [31:0]   _zz_1837;
  wire       [31:0]   _zz_1838;
  wire       [31:0]   _zz_1839;
  wire       [31:0]   _zz_1840;
  wire       [31:0]   _zz_1841;
  wire       [31:0]   _zz_1842;
  wire       [31:0]   _zz_1843;
  wire       [31:0]   _zz_1844;
  wire       [31:0]   _zz_1845;
  wire       [31:0]   _zz_1846;
  wire       [31:0]   _zz_1847;
  wire       [31:0]   _zz_1848;
  wire       [31:0]   _zz_1849;
  wire       [31:0]   _zz_1850;
  wire       [31:0]   _zz_1851;
  wire       [31:0]   _zz_1852;
  wire       [31:0]   _zz_1853;
  wire       [31:0]   _zz_1854;
  wire       [31:0]   _zz_1855;
  wire       [31:0]   _zz_1856;
  wire       [31:0]   _zz_1857;
  wire       [31:0]   _zz_1858;
  wire       [31:0]   _zz_1859;
  wire       [31:0]   _zz_1860;
  wire       [31:0]   _zz_1861;
  wire       [31:0]   _zz_1862;
  wire       [31:0]   _zz_1863;
  wire       [31:0]   _zz_1864;
  wire       [31:0]   _zz_1865;
  wire       [31:0]   _zz_1866;
  wire       [31:0]   _zz_1867;
  wire       [31:0]   _zz_1868;
  wire       [31:0]   _zz_1869;
  wire       [31:0]   _zz_1870;
  wire       [31:0]   _zz_1871;
  wire       [31:0]   _zz_1872;
  wire       [31:0]   _zz_1873;
  wire       [31:0]   _zz_1874;
  wire       [31:0]   _zz_1875;
  wire       [31:0]   _zz_1876;
  wire       [31:0]   _zz_1877;
  wire       [31:0]   _zz_1878;
  wire       [31:0]   _zz_1879;
  wire       [31:0]   _zz_1880;
  wire       [31:0]   _zz_1881;
  wire       [31:0]   _zz_1882;
  wire       [31:0]   _zz_1883;
  wire       [31:0]   _zz_1884;
  wire       [31:0]   _zz_1885;
  wire       [31:0]   _zz_1886;
  wire       [31:0]   _zz_1887;
  wire       [31:0]   _zz_1888;
  wire       [31:0]   _zz_1889;
  wire       [31:0]   _zz_1890;
  wire       [31:0]   _zz_1891;
  wire       [31:0]   _zz_1892;
  wire       [31:0]   _zz_1893;
  wire       [31:0]   _zz_1894;
  wire       [31:0]   _zz_1895;
  wire       [31:0]   _zz_1896;
  wire       [31:0]   _zz_1897;
  wire       [31:0]   _zz_1898;
  wire       [31:0]   _zz_1899;
  wire       [31:0]   _zz_1900;
  wire       [31:0]   _zz_1901;
  wire       [31:0]   _zz_1902;
  wire       [31:0]   _zz_1903;
  wire       [31:0]   _zz_1904;
  wire       [31:0]   _zz_1905;
  wire       [31:0]   _zz_1906;
  wire       [31:0]   _zz_1907;
  wire       [31:0]   _zz_1908;
  wire       [31:0]   _zz_1909;
  wire       [31:0]   _zz_1910;
  wire       [31:0]   _zz_1911;
  wire       [31:0]   _zz_1912;
  wire       [31:0]   _zz_1913;
  wire       [31:0]   _zz_1914;
  wire       [31:0]   _zz_1915;
  wire       [31:0]   _zz_1916;
  wire       [31:0]   _zz_1917;
  wire       [31:0]   _zz_1918;
  wire       [31:0]   _zz_1919;
  wire       [31:0]   _zz_1920;
  wire       [31:0]   _zz_1921;
  wire       [31:0]   _zz_1922;
  wire       [31:0]   _zz_1923;
  wire       [31:0]   _zz_1924;
  wire       [31:0]   _zz_1925;
  wire       [31:0]   _zz_1926;
  wire       [31:0]   _zz_1927;
  wire       [31:0]   _zz_1928;
  wire       [31:0]   _zz_1929;
  wire       [31:0]   _zz_1930;
  wire       [31:0]   _zz_1931;
  wire       [31:0]   _zz_1932;
  wire       [31:0]   _zz_1933;
  wire       [31:0]   _zz_1934;
  wire       [31:0]   _zz_1935;
  wire       [31:0]   _zz_1936;
  wire       [31:0]   _zz_1937;
  wire       [31:0]   _zz_1938;
  wire       [31:0]   _zz_1939;
  wire       [31:0]   _zz_1940;
  wire       [31:0]   _zz_1941;
  wire       [31:0]   _zz_1942;
  wire       [31:0]   _zz_1943;
  wire       [31:0]   _zz_1944;
  wire       [31:0]   _zz_1945;
  wire       [31:0]   _zz_1946;
  wire       [31:0]   _zz_1947;
  wire       [31:0]   _zz_1948;
  wire       [31:0]   _zz_1949;
  wire       [31:0]   _zz_1950;
  wire       [31:0]   _zz_1951;
  wire       [31:0]   _zz_1952;
  wire       [31:0]   _zz_1953;
  wire       [31:0]   _zz_1954;
  wire       [31:0]   _zz_1955;
  wire       [31:0]   _zz_1956;
  wire       [31:0]   _zz_1957;
  wire       [31:0]   _zz_1958;
  wire       [31:0]   _zz_1959;
  wire       [31:0]   _zz_1960;
  wire       [31:0]   _zz_1961;
  wire       [31:0]   _zz_1962;
  wire       [31:0]   _zz_1963;
  wire       [31:0]   _zz_1964;
  wire       [31:0]   _zz_1965;
  wire       [31:0]   _zz_1966;
  wire       [31:0]   _zz_1967;
  wire       [31:0]   _zz_1968;
  wire       [31:0]   _zz_1969;
  wire       [31:0]   _zz_1970;
  wire       [31:0]   _zz_1971;
  wire       [31:0]   _zz_1972;
  wire       [31:0]   _zz_1973;
  wire       [31:0]   _zz_1974;
  wire       [31:0]   _zz_1975;
  wire       [31:0]   _zz_1976;
  wire       [31:0]   _zz_1977;
  wire       [31:0]   _zz_1978;
  wire       [31:0]   _zz_1979;
  wire       [31:0]   _zz_1980;
  wire       [31:0]   _zz_1981;
  wire       [31:0]   _zz_1982;
  wire       [31:0]   _zz_1983;
  wire       [31:0]   _zz_1984;
  wire       [31:0]   _zz_1985;
  wire       [31:0]   _zz_1986;
  wire       [31:0]   _zz_1987;
  wire       [31:0]   _zz_1988;
  wire       [31:0]   _zz_1989;
  wire       [31:0]   _zz_1990;
  wire       [31:0]   _zz_1991;
  wire       [31:0]   _zz_1992;
  wire       [31:0]   _zz_1993;
  wire       [31:0]   _zz_1994;
  wire       [31:0]   _zz_1995;
  wire       [31:0]   _zz_1996;
  wire       [31:0]   _zz_1997;
  wire       [31:0]   _zz_1998;
  wire       [31:0]   _zz_1999;
  wire       [31:0]   _zz_2000;
  wire       [31:0]   _zz_2001;
  wire       [31:0]   _zz_2002;
  wire       [31:0]   _zz_2003;
  wire       [31:0]   _zz_2004;
  wire       [31:0]   _zz_2005;
  wire       [31:0]   _zz_2006;
  wire       [31:0]   _zz_2007;
  wire       [31:0]   _zz_2008;
  wire       [31:0]   _zz_2009;
  wire       [31:0]   _zz_2010;
  wire       [31:0]   _zz_2011;
  wire       [31:0]   _zz_2012;
  wire       [31:0]   _zz_2013;
  wire       [31:0]   _zz_2014;
  wire       [31:0]   _zz_2015;
  wire       [31:0]   _zz_2016;
  wire       [31:0]   _zz_2017;
  wire       [31:0]   _zz_2018;
  wire       [31:0]   _zz_2019;
  wire       [31:0]   _zz_2020;
  wire       [31:0]   _zz_2021;
  wire       [31:0]   _zz_2022;
  wire       [31:0]   _zz_2023;
  wire       [31:0]   _zz_2024;
  wire       [31:0]   _zz_2025;
  wire       [31:0]   _zz_2026;
  wire       [31:0]   _zz_2027;
  wire       [31:0]   _zz_2028;
  wire       [31:0]   _zz_2029;
  wire       [31:0]   _zz_2030;
  wire       [31:0]   _zz_2031;
  wire       [31:0]   _zz_2032;
  wire       [31:0]   _zz_2033;
  wire       [31:0]   _zz_2034;
  wire       [31:0]   _zz_2035;
  wire       [31:0]   _zz_2036;
  wire       [31:0]   _zz_2037;
  wire       [31:0]   _zz_2038;
  wire       [31:0]   _zz_2039;
  wire       [31:0]   _zz_2040;
  wire       [31:0]   _zz_2041;
  wire       [31:0]   _zz_2042;
  wire       [31:0]   _zz_2043;
  wire       [31:0]   _zz_2044;
  wire       [31:0]   _zz_2045;
  wire       [31:0]   _zz_2046;
  wire       [31:0]   _zz_2047;
  wire       [31:0]   _zz_2048;
  wire       [31:0]   _zz_2049;
  wire       [31:0]   _zz_2050;
  wire       [31:0]   _zz_2051;
  wire       [31:0]   _zz_2052;
  wire       [31:0]   _zz_2053;
  wire       [31:0]   _zz_2054;
  wire       [31:0]   _zz_2055;
  wire       [31:0]   _zz_2056;
  wire       [31:0]   _zz_2057;
  wire       [31:0]   _zz_2058;
  wire       [31:0]   _zz_2059;
  wire       [31:0]   _zz_2060;
  wire       [31:0]   _zz_2061;
  wire       [31:0]   _zz_2062;
  wire       [31:0]   _zz_2063;
  wire       [31:0]   _zz_2064;
  wire       [31:0]   _zz_2065;
  wire       [31:0]   _zz_2066;
  wire       [31:0]   _zz_2067;
  wire       [31:0]   _zz_2068;
  wire       [31:0]   _zz_2069;
  wire       [31:0]   _zz_2070;
  wire       [31:0]   _zz_2071;
  wire       [31:0]   _zz_2072;
  wire       [31:0]   _zz_2073;
  wire       [31:0]   _zz_2074;
  wire       [31:0]   _zz_2075;
  wire       [31:0]   _zz_2076;
  wire       [31:0]   _zz_2077;
  wire       [31:0]   _zz_2078;
  wire       [31:0]   _zz_2079;
  wire       [31:0]   _zz_2080;
  wire       [31:0]   _zz_2081;
  wire       [31:0]   _zz_2082;
  wire       [31:0]   _zz_2083;
  wire       [31:0]   _zz_2084;
  wire       [31:0]   _zz_2085;
  wire       [31:0]   _zz_2086;
  wire       [31:0]   _zz_2087;
  wire       [31:0]   _zz_2088;
  wire       [31:0]   _zz_2089;
  wire       [31:0]   _zz_2090;
  wire       [31:0]   _zz_2091;
  wire       [31:0]   _zz_2092;
  wire       [31:0]   _zz_2093;
  wire       [31:0]   _zz_2094;
  wire       [31:0]   _zz_2095;
  wire       [31:0]   _zz_2096;
  wire       [31:0]   _zz_2097;
  wire       [31:0]   _zz_2098;
  wire       [31:0]   _zz_2099;
  wire       [31:0]   _zz_2100;
  wire       [31:0]   _zz_2101;
  wire       [31:0]   _zz_2102;
  wire       [31:0]   _zz_2103;
  wire       [31:0]   _zz_2104;
  wire       [31:0]   _zz_2105;
  wire       [31:0]   _zz_2106;
  wire       [31:0]   _zz_2107;
  wire       [31:0]   _zz_2108;
  wire       [31:0]   _zz_2109;
  wire       [31:0]   _zz_2110;
  wire       [31:0]   _zz_2111;
  wire       [31:0]   _zz_2112;
  wire       [31:0]   _zz_2113;
  wire       [31:0]   _zz_2114;
  wire       [31:0]   _zz_2115;
  wire       [31:0]   _zz_2116;
  wire       [31:0]   _zz_2117;
  wire       [31:0]   _zz_2118;
  wire       [31:0]   _zz_2119;
  wire       [31:0]   _zz_2120;
  wire       [31:0]   _zz_2121;
  wire       [31:0]   _zz_2122;
  wire       [31:0]   _zz_2123;
  wire       [31:0]   _zz_2124;
  wire       [31:0]   _zz_2125;
  wire       [31:0]   _zz_2126;
  wire       [31:0]   _zz_2127;
  wire       [31:0]   _zz_2128;
  wire       [31:0]   _zz_2129;
  wire       [31:0]   _zz_2130;
  wire       [31:0]   _zz_2131;
  wire       [31:0]   _zz_2132;
  wire       [31:0]   _zz_2133;
  wire       [31:0]   _zz_2134;
  wire       [31:0]   _zz_2135;
  wire       [31:0]   _zz_2136;
  wire       [31:0]   _zz_2137;
  wire       [31:0]   _zz_2138;
  wire       [31:0]   _zz_2139;
  wire       [31:0]   _zz_2140;
  wire       [31:0]   _zz_2141;
  wire       [31:0]   _zz_2142;
  wire       [31:0]   _zz_2143;
  wire       [31:0]   _zz_2144;
  wire       [31:0]   _zz_2145;
  wire       [31:0]   _zz_2146;
  wire       [31:0]   _zz_2147;
  wire       [31:0]   _zz_2148;
  wire       [31:0]   _zz_2149;
  wire       [31:0]   _zz_2150;
  wire       [31:0]   _zz_2151;
  wire       [31:0]   _zz_2152;
  wire       [31:0]   _zz_2153;
  wire       [31:0]   _zz_2154;
  wire       [31:0]   _zz_2155;
  wire       [31:0]   _zz_2156;
  wire       [31:0]   _zz_2157;
  wire       [31:0]   _zz_2158;
  wire       [31:0]   _zz_2159;
  wire       [31:0]   _zz_2160;
  wire       [31:0]   _zz_2161;
  wire       [31:0]   _zz_2162;
  wire       [31:0]   _zz_2163;
  wire       [31:0]   _zz_2164;
  wire       [31:0]   _zz_2165;
  wire       [31:0]   _zz_2166;
  wire       [31:0]   _zz_2167;
  wire       [31:0]   _zz_2168;
  wire       [31:0]   _zz_2169;
  wire       [31:0]   _zz_2170;
  wire       [31:0]   _zz_2171;
  wire       [31:0]   _zz_2172;
  wire       [31:0]   _zz_2173;
  wire       [31:0]   _zz_2174;
  wire       [31:0]   _zz_2175;
  wire       [31:0]   _zz_2176;
  wire       [31:0]   _zz_2177;
  wire       [31:0]   _zz_2178;
  wire       [31:0]   _zz_2179;
  wire       [31:0]   _zz_2180;
  wire       [31:0]   _zz_2181;
  wire       [31:0]   _zz_2182;
  wire       [31:0]   _zz_2183;
  wire       [31:0]   _zz_2184;
  wire       [31:0]   _zz_2185;
  wire       [31:0]   _zz_2186;
  wire       [31:0]   _zz_2187;
  wire       [31:0]   _zz_2188;
  wire       [31:0]   _zz_2189;
  wire       [31:0]   _zz_2190;
  wire       [31:0]   _zz_2191;
  wire       [31:0]   _zz_2192;
  wire       [31:0]   _zz_2193;
  wire       [31:0]   _zz_2194;
  wire       [31:0]   _zz_2195;
  wire       [31:0]   _zz_2196;
  wire       [31:0]   _zz_2197;
  wire       [31:0]   _zz_2198;
  wire       [31:0]   _zz_2199;
  wire       [31:0]   _zz_2200;
  wire       [31:0]   _zz_2201;
  wire       [31:0]   _zz_2202;
  wire       [31:0]   _zz_2203;
  wire       [31:0]   _zz_2204;
  wire       [31:0]   _zz_2205;
  wire       [31:0]   _zz_2206;
  wire       [31:0]   _zz_2207;
  wire       [31:0]   _zz_2208;
  wire       [31:0]   _zz_2209;
  wire       [31:0]   _zz_2210;
  wire       [31:0]   _zz_2211;
  wire       [31:0]   _zz_2212;
  wire       [31:0]   _zz_2213;
  wire       [31:0]   _zz_2214;
  wire       [31:0]   _zz_2215;
  wire       [31:0]   _zz_2216;
  wire       [31:0]   _zz_2217;
  wire       [31:0]   _zz_2218;
  wire       [31:0]   _zz_2219;
  wire       [31:0]   _zz_2220;
  wire       [31:0]   _zz_2221;
  wire       [31:0]   _zz_2222;
  wire       [31:0]   _zz_2223;
  wire       [31:0]   _zz_2224;
  wire       [31:0]   _zz_2225;
  wire       [31:0]   _zz_2226;
  wire       [31:0]   _zz_2227;
  wire       [31:0]   _zz_2228;
  wire       [31:0]   _zz_2229;
  wire       [31:0]   _zz_2230;
  wire       [31:0]   _zz_2231;
  wire       [31:0]   _zz_2232;
  wire       [31:0]   _zz_2233;
  wire       [31:0]   _zz_2234;
  wire       [31:0]   _zz_2235;
  wire       [31:0]   _zz_2236;
  wire       [31:0]   _zz_2237;
  wire       [31:0]   _zz_2238;
  wire       [31:0]   _zz_2239;
  wire       [31:0]   _zz_2240;
  wire       [31:0]   _zz_2241;
  wire       [31:0]   _zz_2242;
  wire       [31:0]   _zz_2243;
  wire       [31:0]   _zz_2244;
  wire       [31:0]   _zz_2245;
  wire       [31:0]   _zz_2246;
  wire       [31:0]   _zz_2247;
  wire       [31:0]   _zz_2248;
  wire       [31:0]   _zz_2249;
  wire       [31:0]   _zz_2250;
  wire       [31:0]   _zz_2251;
  wire       [31:0]   _zz_2252;
  wire       [31:0]   _zz_2253;
  wire       [31:0]   _zz_2254;
  wire       [31:0]   _zz_2255;
  wire       [31:0]   _zz_2256;
  wire       [31:0]   _zz_2257;
  wire       [31:0]   _zz_2258;
  wire       [31:0]   _zz_2259;
  wire       [31:0]   _zz_2260;
  wire       [31:0]   _zz_2261;
  wire       [31:0]   _zz_2262;
  wire       [31:0]   _zz_2263;
  wire       [31:0]   _zz_2264;
  wire       [31:0]   _zz_2265;
  wire       [31:0]   _zz_2266;
  wire       [31:0]   _zz_2267;
  wire       [31:0]   _zz_2268;
  wire       [31:0]   _zz_2269;
  wire       [31:0]   _zz_2270;
  wire       [31:0]   _zz_2271;
  wire       [31:0]   _zz_2272;
  wire       [31:0]   _zz_2273;
  wire       [31:0]   _zz_2274;
  wire       [31:0]   _zz_2275;
  wire       [31:0]   _zz_2276;
  wire       [31:0]   _zz_2277;
  wire       [31:0]   _zz_2278;
  wire       [31:0]   _zz_2279;
  wire       [31:0]   _zz_2280;
  wire       [31:0]   _zz_2281;
  wire       [31:0]   _zz_2282;
  wire       [31:0]   _zz_2283;
  wire       [31:0]   _zz_2284;
  wire       [31:0]   _zz_2285;
  wire       [31:0]   _zz_2286;
  wire       [31:0]   _zz_2287;
  wire       [31:0]   _zz_2288;
  wire       [31:0]   _zz_2289;
  wire       [31:0]   _zz_2290;
  wire       [31:0]   _zz_2291;
  wire       [31:0]   _zz_2292;
  wire       [31:0]   _zz_2293;
  wire       [31:0]   _zz_2294;
  wire       [31:0]   _zz_2295;
  wire       [31:0]   _zz_2296;
  wire       [31:0]   _zz_2297;
  wire       [31:0]   _zz_2298;
  wire       [31:0]   _zz_2299;
  wire       [31:0]   _zz_2300;
  wire       [31:0]   _zz_2301;
  wire       [31:0]   _zz_2302;
  wire       [31:0]   _zz_2303;
  wire       [31:0]   _zz_2304;
  wire       [31:0]   _zz_2305;
  wire       [31:0]   _zz_2306;
  wire       [31:0]   _zz_2307;
  wire       [31:0]   _zz_2308;
  wire       [31:0]   _zz_2309;
  wire       [31:0]   _zz_2310;
  wire       [31:0]   _zz_2311;
  wire       [31:0]   _zz_2312;
  wire       [31:0]   _zz_2313;
  wire       [31:0]   _zz_2314;
  wire       [31:0]   _zz_2315;
  wire       [31:0]   _zz_2316;
  wire       [31:0]   _zz_2317;
  wire       [31:0]   _zz_2318;
  wire       [31:0]   _zz_2319;
  wire       [31:0]   _zz_2320;
  wire       [31:0]   _zz_2321;
  wire       [31:0]   _zz_2322;
  wire       [31:0]   _zz_2323;
  wire       [31:0]   _zz_2324;
  wire       [31:0]   _zz_2325;
  wire       [31:0]   _zz_2326;
  wire       [31:0]   _zz_2327;
  wire       [31:0]   _zz_2328;
  wire       [31:0]   _zz_2329;
  wire       [31:0]   _zz_2330;
  wire       [31:0]   _zz_2331;
  wire       [31:0]   _zz_2332;
  wire       [31:0]   _zz_2333;
  wire       [31:0]   _zz_2334;
  wire       [31:0]   _zz_2335;
  wire       [31:0]   _zz_2336;
  wire       [31:0]   _zz_2337;
  wire       [31:0]   _zz_2338;
  wire       [31:0]   _zz_2339;
  wire       [31:0]   _zz_2340;
  wire       [31:0]   _zz_2341;
  wire       [31:0]   _zz_2342;
  wire       [31:0]   _zz_2343;
  wire       [31:0]   _zz_2344;
  wire       [31:0]   _zz_2345;
  wire       [31:0]   _zz_2346;
  wire       [31:0]   _zz_2347;
  wire       [31:0]   _zz_2348;
  wire       [31:0]   _zz_2349;
  wire       [31:0]   _zz_2350;
  wire       [31:0]   _zz_2351;
  wire       [31:0]   _zz_2352;
  wire       [31:0]   _zz_2353;
  wire       [31:0]   _zz_2354;
  wire       [31:0]   _zz_2355;
  wire       [31:0]   _zz_2356;
  wire       [31:0]   _zz_2357;
  wire       [31:0]   _zz_2358;
  wire       [31:0]   _zz_2359;
  wire       [31:0]   _zz_2360;
  wire       [31:0]   _zz_2361;
  wire       [31:0]   _zz_2362;
  wire       [31:0]   _zz_2363;
  wire       [31:0]   _zz_2364;
  wire       [31:0]   _zz_2365;
  wire       [31:0]   _zz_2366;
  wire       [31:0]   _zz_2367;
  wire       [31:0]   _zz_2368;
  wire       [31:0]   _zz_2369;
  wire       [31:0]   _zz_2370;
  wire       [31:0]   _zz_2371;
  wire       [31:0]   _zz_2372;
  wire       [31:0]   _zz_2373;
  wire       [31:0]   _zz_2374;
  wire       [31:0]   _zz_2375;
  wire       [31:0]   _zz_2376;
  wire       [31:0]   _zz_2377;
  wire       [31:0]   _zz_2378;
  wire       [31:0]   _zz_2379;
  wire       [31:0]   _zz_2380;
  wire       [31:0]   _zz_2381;
  wire       [31:0]   _zz_2382;
  wire       [31:0]   _zz_2383;
  wire       [31:0]   _zz_2384;
  wire       [31:0]   _zz_2385;
  wire       [31:0]   _zz_2386;
  wire       [31:0]   _zz_2387;
  wire       [31:0]   _zz_2388;
  wire       [31:0]   _zz_2389;
  wire       [31:0]   _zz_2390;
  wire       [31:0]   _zz_2391;
  wire       [31:0]   _zz_2392;
  wire       [31:0]   _zz_2393;
  wire       [31:0]   _zz_2394;
  wire       [31:0]   _zz_2395;
  wire       [31:0]   _zz_2396;
  wire       [31:0]   _zz_2397;
  wire       [31:0]   _zz_2398;
  wire       [31:0]   _zz_2399;
  wire       [31:0]   _zz_2400;
  wire       [31:0]   _zz_2401;
  wire       [31:0]   _zz_2402;
  wire       [31:0]   _zz_2403;
  wire       [31:0]   _zz_2404;
  wire       [31:0]   _zz_2405;
  wire       [31:0]   _zz_2406;
  wire       [31:0]   _zz_2407;
  wire       [31:0]   _zz_2408;
  wire       [31:0]   _zz_2409;
  wire       [31:0]   _zz_2410;
  wire       [31:0]   _zz_2411;
  wire       [31:0]   _zz_2412;
  wire       [31:0]   _zz_2413;
  wire       [31:0]   _zz_2414;
  wire       [31:0]   _zz_2415;
  wire       [31:0]   _zz_2416;
  wire       [31:0]   _zz_2417;
  wire       [31:0]   _zz_2418;
  wire       [31:0]   _zz_2419;
  wire       [31:0]   _zz_2420;
  wire       [31:0]   _zz_2421;
  wire       [31:0]   _zz_2422;
  wire       [31:0]   _zz_2423;
  wire       [31:0]   _zz_2424;
  wire       [31:0]   _zz_2425;
  wire       [31:0]   _zz_2426;
  wire       [31:0]   _zz_2427;
  wire       [31:0]   _zz_2428;
  wire       [31:0]   _zz_2429;
  wire       [31:0]   _zz_2430;
  wire       [31:0]   _zz_2431;
  wire       [31:0]   _zz_2432;
  wire       [31:0]   _zz_2433;
  wire       [31:0]   _zz_2434;
  wire       [31:0]   _zz_2435;
  wire       [31:0]   _zz_2436;
  wire       [31:0]   _zz_2437;
  wire       [31:0]   _zz_2438;
  wire       [31:0]   _zz_2439;
  wire       [31:0]   _zz_2440;
  wire       [31:0]   _zz_2441;
  wire       [31:0]   _zz_2442;
  wire       [31:0]   _zz_2443;
  wire       [31:0]   _zz_2444;
  wire       [31:0]   _zz_2445;
  wire       [31:0]   _zz_2446;
  wire       [31:0]   _zz_2447;
  wire       [31:0]   _zz_2448;
  wire       [31:0]   _zz_2449;
  wire       [31:0]   _zz_2450;
  wire       [31:0]   _zz_2451;
  wire       [31:0]   _zz_2452;
  wire       [31:0]   _zz_2453;
  wire       [31:0]   _zz_2454;
  wire       [31:0]   _zz_2455;
  wire       [31:0]   _zz_2456;
  wire       [31:0]   _zz_2457;
  wire       [31:0]   _zz_2458;
  wire       [31:0]   _zz_2459;
  wire       [31:0]   _zz_2460;
  wire       [31:0]   _zz_2461;
  wire       [31:0]   _zz_2462;
  wire       [31:0]   _zz_2463;
  wire       [31:0]   _zz_2464;
  wire       [31:0]   _zz_2465;
  wire       [31:0]   _zz_2466;
  wire       [31:0]   _zz_2467;
  wire       [31:0]   _zz_2468;
  wire       [31:0]   _zz_2469;
  wire       [31:0]   _zz_2470;
  wire       [31:0]   _zz_2471;
  wire       [31:0]   _zz_2472;
  wire       [31:0]   _zz_2473;
  wire       [31:0]   _zz_2474;
  wire       [31:0]   _zz_2475;
  wire       [31:0]   _zz_2476;
  wire       [31:0]   _zz_2477;
  wire       [31:0]   _zz_2478;
  wire       [31:0]   _zz_2479;
  wire       [31:0]   _zz_2480;
  wire       [31:0]   _zz_2481;
  wire       [31:0]   _zz_2482;
  wire       [31:0]   _zz_2483;
  wire       [31:0]   _zz_2484;
  wire       [31:0]   _zz_2485;
  wire       [31:0]   _zz_2486;
  wire       [31:0]   _zz_2487;
  wire       [31:0]   _zz_2488;
  wire       [31:0]   _zz_2489;
  wire       [31:0]   _zz_2490;
  wire       [31:0]   _zz_2491;
  wire       [31:0]   _zz_2492;
  wire       [31:0]   _zz_2493;
  wire       [31:0]   _zz_2494;
  wire       [31:0]   _zz_2495;
  wire       [31:0]   _zz_2496;
  wire       [31:0]   _zz_2497;
  wire       [31:0]   _zz_2498;
  wire       [31:0]   _zz_2499;
  wire       [31:0]   _zz_2500;
  wire       [31:0]   _zz_2501;
  wire       [31:0]   _zz_2502;
  wire       [31:0]   _zz_2503;
  wire       [31:0]   _zz_2504;
  wire       [31:0]   _zz_2505;
  wire       [31:0]   _zz_2506;
  wire       [31:0]   _zz_2507;
  wire       [31:0]   _zz_2508;
  wire       [31:0]   _zz_2509;
  wire       [31:0]   _zz_2510;
  wire       [31:0]   _zz_2511;
  wire       [31:0]   _zz_2512;
  wire       [31:0]   _zz_2513;
  wire       [31:0]   _zz_2514;
  wire       [31:0]   _zz_2515;
  wire       [31:0]   _zz_2516;
  wire       [31:0]   _zz_2517;
  wire       [31:0]   _zz_2518;
  wire       [31:0]   _zz_2519;
  wire       [31:0]   _zz_2520;
  wire       [31:0]   _zz_2521;
  wire       [31:0]   _zz_2522;
  wire       [31:0]   _zz_2523;
  wire       [31:0]   _zz_2524;
  wire       [31:0]   _zz_2525;
  wire       [31:0]   _zz_2526;
  wire       [31:0]   _zz_2527;
  wire       [31:0]   _zz_2528;
  wire       [31:0]   _zz_2529;
  wire       [31:0]   _zz_2530;
  wire       [31:0]   _zz_2531;
  wire       [31:0]   _zz_2532;
  wire       [31:0]   _zz_2533;
  wire       [31:0]   _zz_2534;
  wire       [31:0]   _zz_2535;
  wire       [31:0]   _zz_2536;
  wire       [31:0]   _zz_2537;
  wire       [31:0]   _zz_2538;
  wire       [31:0]   _zz_2539;
  wire       [31:0]   _zz_2540;
  wire       [31:0]   _zz_2541;
  wire       [31:0]   _zz_2542;
  wire       [31:0]   _zz_2543;
  wire       [31:0]   _zz_2544;
  wire       [31:0]   _zz_2545;
  wire       [31:0]   _zz_2546;
  wire       [31:0]   _zz_2547;
  wire       [31:0]   _zz_2548;
  wire       [31:0]   _zz_2549;
  wire       [31:0]   _zz_2550;
  wire       [31:0]   _zz_2551;
  wire       [31:0]   _zz_2552;
  wire       [31:0]   _zz_2553;
  wire       [31:0]   _zz_2554;
  wire       [31:0]   _zz_2555;
  wire       [31:0]   _zz_2556;
  wire       [31:0]   _zz_2557;
  wire       [31:0]   _zz_2558;
  wire       [31:0]   _zz_2559;
  wire       [31:0]   _zz_2560;
  wire       [31:0]   _zz_2561;
  wire       [31:0]   _zz_2562;
  wire       [31:0]   _zz_2563;
  wire       [31:0]   _zz_2564;
  wire       [31:0]   _zz_2565;
  wire       [31:0]   _zz_2566;
  wire       [31:0]   _zz_2567;
  wire       [31:0]   _zz_2568;
  wire       [31:0]   _zz_2569;
  wire       [31:0]   _zz_2570;
  wire       [31:0]   _zz_2571;
  wire       [31:0]   _zz_2572;
  wire       [31:0]   _zz_2573;
  wire       [31:0]   _zz_2574;
  wire       [31:0]   _zz_2575;
  wire       [31:0]   _zz_2576;
  wire       [31:0]   _zz_2577;
  wire       [31:0]   _zz_2578;
  wire       [31:0]   _zz_2579;
  wire       [31:0]   _zz_2580;
  wire       [31:0]   _zz_2581;
  wire       [31:0]   _zz_2582;
  wire       [31:0]   _zz_2583;
  wire       [31:0]   _zz_2584;
  wire       [31:0]   _zz_2585;
  wire       [31:0]   _zz_2586;
  wire       [31:0]   _zz_2587;
  wire       [31:0]   _zz_2588;
  wire       [31:0]   _zz_2589;
  wire       [31:0]   _zz_2590;
  wire       [31:0]   _zz_2591;
  wire       [31:0]   _zz_2592;
  wire       [31:0]   _zz_2593;
  wire       [31:0]   _zz_2594;
  wire       [31:0]   _zz_2595;
  wire       [31:0]   _zz_2596;
  wire       [31:0]   _zz_2597;
  wire       [31:0]   _zz_2598;
  wire       [31:0]   _zz_2599;
  wire       [31:0]   _zz_2600;
  wire       [31:0]   _zz_2601;
  wire       [31:0]   _zz_2602;
  wire       [31:0]   _zz_2603;
  wire       [31:0]   _zz_2604;
  wire       [31:0]   _zz_2605;
  wire       [31:0]   _zz_2606;
  wire       [31:0]   _zz_2607;
  wire       [31:0]   _zz_2608;
  wire       [31:0]   _zz_2609;
  wire       [31:0]   _zz_2610;
  wire       [31:0]   _zz_2611;
  wire       [31:0]   _zz_2612;
  wire       [31:0]   _zz_2613;
  wire       [31:0]   _zz_2614;
  wire       [31:0]   _zz_2615;
  wire       [31:0]   _zz_2616;
  wire       [31:0]   _zz_2617;
  wire       [31:0]   _zz_2618;
  wire       [31:0]   _zz_2619;
  wire       [31:0]   _zz_2620;
  wire       [31:0]   _zz_2621;
  wire       [31:0]   _zz_2622;
  wire       [31:0]   _zz_2623;
  wire       [31:0]   _zz_2624;
  wire       [31:0]   _zz_2625;
  wire       [31:0]   _zz_2626;
  wire       [31:0]   _zz_2627;
  wire       [31:0]   _zz_2628;
  wire       [31:0]   _zz_2629;
  wire       [31:0]   _zz_2630;
  wire       [31:0]   _zz_2631;
  wire       [31:0]   _zz_2632;
  wire       [31:0]   _zz_2633;
  wire       [31:0]   _zz_2634;
  wire       [31:0]   _zz_2635;
  wire       [31:0]   _zz_2636;
  wire       [31:0]   _zz_2637;
  wire       [31:0]   _zz_2638;
  wire       [31:0]   _zz_2639;
  wire       [31:0]   _zz_2640;
  wire       [31:0]   _zz_2641;
  wire       [31:0]   _zz_2642;
  wire       [31:0]   _zz_2643;
  wire       [31:0]   _zz_2644;
  wire       [31:0]   _zz_2645;
  wire       [31:0]   _zz_2646;
  wire       [31:0]   _zz_2647;
  wire       [31:0]   _zz_2648;
  wire       [31:0]   _zz_2649;
  wire       [31:0]   _zz_2650;
  wire       [31:0]   _zz_2651;
  wire       [31:0]   _zz_2652;
  wire       [31:0]   _zz_2653;
  wire       [31:0]   _zz_2654;
  wire       [31:0]   _zz_2655;
  wire       [31:0]   _zz_2656;
  wire       [31:0]   _zz_2657;
  wire       [31:0]   _zz_2658;
  wire       [31:0]   _zz_2659;
  wire       [31:0]   _zz_2660;
  wire       [31:0]   _zz_2661;
  wire       [31:0]   _zz_2662;
  wire       [31:0]   _zz_2663;
  wire       [31:0]   _zz_2664;
  wire       [31:0]   _zz_2665;
  wire       [31:0]   _zz_2666;
  wire       [31:0]   _zz_2667;
  wire       [31:0]   _zz_2668;
  wire       [31:0]   _zz_2669;
  wire       [31:0]   _zz_2670;
  wire       [31:0]   _zz_2671;
  wire       [31:0]   _zz_2672;
  wire       [31:0]   _zz_2673;
  wire       [31:0]   _zz_2674;
  wire       [31:0]   _zz_2675;
  wire       [31:0]   _zz_2676;
  wire       [31:0]   _zz_2677;
  wire       [31:0]   _zz_2678;
  wire       [31:0]   _zz_2679;
  wire       [31:0]   _zz_2680;
  wire       [31:0]   _zz_2681;
  wire       [31:0]   _zz_2682;
  wire       [31:0]   _zz_2683;
  wire       [31:0]   _zz_2684;
  wire       [31:0]   _zz_2685;
  wire       [31:0]   _zz_2686;
  wire       [31:0]   _zz_2687;
  wire       [31:0]   _zz_2688;
  wire       [15:0]   fixTo_dout;
  wire       [15:0]   fixTo_1_dout;
  wire       [15:0]   fixTo_2_dout;
  wire       [15:0]   fixTo_3_dout;
  wire       [15:0]   fixTo_4_dout;
  wire       [15:0]   fixTo_5_dout;
  wire       [15:0]   fixTo_6_dout;
  wire       [15:0]   fixTo_7_dout;
  wire       [15:0]   fixTo_8_dout;
  wire       [15:0]   fixTo_9_dout;
  wire       [15:0]   fixTo_10_dout;
  wire       [15:0]   fixTo_11_dout;
  wire       [15:0]   fixTo_12_dout;
  wire       [15:0]   fixTo_13_dout;
  wire       [15:0]   fixTo_14_dout;
  wire       [15:0]   fixTo_15_dout;
  wire       [15:0]   fixTo_16_dout;
  wire       [15:0]   fixTo_17_dout;
  wire       [15:0]   fixTo_18_dout;
  wire       [15:0]   fixTo_19_dout;
  wire       [15:0]   fixTo_20_dout;
  wire       [15:0]   fixTo_21_dout;
  wire       [15:0]   fixTo_22_dout;
  wire       [15:0]   fixTo_23_dout;
  wire       [15:0]   fixTo_24_dout;
  wire       [15:0]   fixTo_25_dout;
  wire       [15:0]   fixTo_26_dout;
  wire       [15:0]   fixTo_27_dout;
  wire       [15:0]   fixTo_28_dout;
  wire       [15:0]   fixTo_29_dout;
  wire       [15:0]   fixTo_30_dout;
  wire       [15:0]   fixTo_31_dout;
  wire       [15:0]   fixTo_32_dout;
  wire       [15:0]   fixTo_33_dout;
  wire       [15:0]   fixTo_34_dout;
  wire       [15:0]   fixTo_35_dout;
  wire       [15:0]   fixTo_36_dout;
  wire       [15:0]   fixTo_37_dout;
  wire       [15:0]   fixTo_38_dout;
  wire       [15:0]   fixTo_39_dout;
  wire       [15:0]   fixTo_40_dout;
  wire       [15:0]   fixTo_41_dout;
  wire       [15:0]   fixTo_42_dout;
  wire       [15:0]   fixTo_43_dout;
  wire       [15:0]   fixTo_44_dout;
  wire       [15:0]   fixTo_45_dout;
  wire       [15:0]   fixTo_46_dout;
  wire       [15:0]   fixTo_47_dout;
  wire       [15:0]   fixTo_48_dout;
  wire       [15:0]   fixTo_49_dout;
  wire       [15:0]   fixTo_50_dout;
  wire       [15:0]   fixTo_51_dout;
  wire       [15:0]   fixTo_52_dout;
  wire       [15:0]   fixTo_53_dout;
  wire       [15:0]   fixTo_54_dout;
  wire       [15:0]   fixTo_55_dout;
  wire       [15:0]   fixTo_56_dout;
  wire       [15:0]   fixTo_57_dout;
  wire       [15:0]   fixTo_58_dout;
  wire       [15:0]   fixTo_59_dout;
  wire       [15:0]   fixTo_60_dout;
  wire       [15:0]   fixTo_61_dout;
  wire       [15:0]   fixTo_62_dout;
  wire       [15:0]   fixTo_63_dout;
  wire       [15:0]   fixTo_64_dout;
  wire       [15:0]   fixTo_65_dout;
  wire       [15:0]   fixTo_66_dout;
  wire       [15:0]   fixTo_67_dout;
  wire       [15:0]   fixTo_68_dout;
  wire       [15:0]   fixTo_69_dout;
  wire       [15:0]   fixTo_70_dout;
  wire       [15:0]   fixTo_71_dout;
  wire       [15:0]   fixTo_72_dout;
  wire       [15:0]   fixTo_73_dout;
  wire       [15:0]   fixTo_74_dout;
  wire       [15:0]   fixTo_75_dout;
  wire       [15:0]   fixTo_76_dout;
  wire       [15:0]   fixTo_77_dout;
  wire       [15:0]   fixTo_78_dout;
  wire       [15:0]   fixTo_79_dout;
  wire       [15:0]   fixTo_80_dout;
  wire       [15:0]   fixTo_81_dout;
  wire       [15:0]   fixTo_82_dout;
  wire       [15:0]   fixTo_83_dout;
  wire       [15:0]   fixTo_84_dout;
  wire       [15:0]   fixTo_85_dout;
  wire       [15:0]   fixTo_86_dout;
  wire       [15:0]   fixTo_87_dout;
  wire       [15:0]   fixTo_88_dout;
  wire       [15:0]   fixTo_89_dout;
  wire       [15:0]   fixTo_90_dout;
  wire       [15:0]   fixTo_91_dout;
  wire       [15:0]   fixTo_92_dout;
  wire       [15:0]   fixTo_93_dout;
  wire       [15:0]   fixTo_94_dout;
  wire       [15:0]   fixTo_95_dout;
  wire       [15:0]   fixTo_96_dout;
  wire       [15:0]   fixTo_97_dout;
  wire       [15:0]   fixTo_98_dout;
  wire       [15:0]   fixTo_99_dout;
  wire       [15:0]   fixTo_100_dout;
  wire       [15:0]   fixTo_101_dout;
  wire       [15:0]   fixTo_102_dout;
  wire       [15:0]   fixTo_103_dout;
  wire       [15:0]   fixTo_104_dout;
  wire       [15:0]   fixTo_105_dout;
  wire       [15:0]   fixTo_106_dout;
  wire       [15:0]   fixTo_107_dout;
  wire       [15:0]   fixTo_108_dout;
  wire       [15:0]   fixTo_109_dout;
  wire       [15:0]   fixTo_110_dout;
  wire       [15:0]   fixTo_111_dout;
  wire       [15:0]   fixTo_112_dout;
  wire       [15:0]   fixTo_113_dout;
  wire       [15:0]   fixTo_114_dout;
  wire       [15:0]   fixTo_115_dout;
  wire       [15:0]   fixTo_116_dout;
  wire       [15:0]   fixTo_117_dout;
  wire       [15:0]   fixTo_118_dout;
  wire       [15:0]   fixTo_119_dout;
  wire       [15:0]   fixTo_120_dout;
  wire       [15:0]   fixTo_121_dout;
  wire       [15:0]   fixTo_122_dout;
  wire       [15:0]   fixTo_123_dout;
  wire       [15:0]   fixTo_124_dout;
  wire       [15:0]   fixTo_125_dout;
  wire       [15:0]   fixTo_126_dout;
  wire       [15:0]   fixTo_127_dout;
  wire       [15:0]   fixTo_128_dout;
  wire       [15:0]   fixTo_129_dout;
  wire       [15:0]   fixTo_130_dout;
  wire       [15:0]   fixTo_131_dout;
  wire       [15:0]   fixTo_132_dout;
  wire       [15:0]   fixTo_133_dout;
  wire       [15:0]   fixTo_134_dout;
  wire       [15:0]   fixTo_135_dout;
  wire       [15:0]   fixTo_136_dout;
  wire       [15:0]   fixTo_137_dout;
  wire       [15:0]   fixTo_138_dout;
  wire       [15:0]   fixTo_139_dout;
  wire       [15:0]   fixTo_140_dout;
  wire       [15:0]   fixTo_141_dout;
  wire       [15:0]   fixTo_142_dout;
  wire       [15:0]   fixTo_143_dout;
  wire       [15:0]   fixTo_144_dout;
  wire       [15:0]   fixTo_145_dout;
  wire       [15:0]   fixTo_146_dout;
  wire       [15:0]   fixTo_147_dout;
  wire       [15:0]   fixTo_148_dout;
  wire       [15:0]   fixTo_149_dout;
  wire       [15:0]   fixTo_150_dout;
  wire       [15:0]   fixTo_151_dout;
  wire       [15:0]   fixTo_152_dout;
  wire       [15:0]   fixTo_153_dout;
  wire       [15:0]   fixTo_154_dout;
  wire       [15:0]   fixTo_155_dout;
  wire       [15:0]   fixTo_156_dout;
  wire       [15:0]   fixTo_157_dout;
  wire       [15:0]   fixTo_158_dout;
  wire       [15:0]   fixTo_159_dout;
  wire       [15:0]   fixTo_160_dout;
  wire       [15:0]   fixTo_161_dout;
  wire       [15:0]   fixTo_162_dout;
  wire       [15:0]   fixTo_163_dout;
  wire       [15:0]   fixTo_164_dout;
  wire       [15:0]   fixTo_165_dout;
  wire       [15:0]   fixTo_166_dout;
  wire       [15:0]   fixTo_167_dout;
  wire       [15:0]   fixTo_168_dout;
  wire       [15:0]   fixTo_169_dout;
  wire       [15:0]   fixTo_170_dout;
  wire       [15:0]   fixTo_171_dout;
  wire       [15:0]   fixTo_172_dout;
  wire       [15:0]   fixTo_173_dout;
  wire       [15:0]   fixTo_174_dout;
  wire       [15:0]   fixTo_175_dout;
  wire       [15:0]   fixTo_176_dout;
  wire       [15:0]   fixTo_177_dout;
  wire       [15:0]   fixTo_178_dout;
  wire       [15:0]   fixTo_179_dout;
  wire       [15:0]   fixTo_180_dout;
  wire       [15:0]   fixTo_181_dout;
  wire       [15:0]   fixTo_182_dout;
  wire       [15:0]   fixTo_183_dout;
  wire       [15:0]   fixTo_184_dout;
  wire       [15:0]   fixTo_185_dout;
  wire       [15:0]   fixTo_186_dout;
  wire       [15:0]   fixTo_187_dout;
  wire       [15:0]   fixTo_188_dout;
  wire       [15:0]   fixTo_189_dout;
  wire       [15:0]   fixTo_190_dout;
  wire       [15:0]   fixTo_191_dout;
  wire       [15:0]   fixTo_192_dout;
  wire       [15:0]   fixTo_193_dout;
  wire       [15:0]   fixTo_194_dout;
  wire       [15:0]   fixTo_195_dout;
  wire       [15:0]   fixTo_196_dout;
  wire       [15:0]   fixTo_197_dout;
  wire       [15:0]   fixTo_198_dout;
  wire       [15:0]   fixTo_199_dout;
  wire       [15:0]   fixTo_200_dout;
  wire       [15:0]   fixTo_201_dout;
  wire       [15:0]   fixTo_202_dout;
  wire       [15:0]   fixTo_203_dout;
  wire       [15:0]   fixTo_204_dout;
  wire       [15:0]   fixTo_205_dout;
  wire       [15:0]   fixTo_206_dout;
  wire       [15:0]   fixTo_207_dout;
  wire       [15:0]   fixTo_208_dout;
  wire       [15:0]   fixTo_209_dout;
  wire       [15:0]   fixTo_210_dout;
  wire       [15:0]   fixTo_211_dout;
  wire       [15:0]   fixTo_212_dout;
  wire       [15:0]   fixTo_213_dout;
  wire       [15:0]   fixTo_214_dout;
  wire       [15:0]   fixTo_215_dout;
  wire       [15:0]   fixTo_216_dout;
  wire       [15:0]   fixTo_217_dout;
  wire       [15:0]   fixTo_218_dout;
  wire       [15:0]   fixTo_219_dout;
  wire       [15:0]   fixTo_220_dout;
  wire       [15:0]   fixTo_221_dout;
  wire       [15:0]   fixTo_222_dout;
  wire       [15:0]   fixTo_223_dout;
  wire       [15:0]   fixTo_224_dout;
  wire       [15:0]   fixTo_225_dout;
  wire       [15:0]   fixTo_226_dout;
  wire       [15:0]   fixTo_227_dout;
  wire       [15:0]   fixTo_228_dout;
  wire       [15:0]   fixTo_229_dout;
  wire       [15:0]   fixTo_230_dout;
  wire       [15:0]   fixTo_231_dout;
  wire       [15:0]   fixTo_232_dout;
  wire       [15:0]   fixTo_233_dout;
  wire       [15:0]   fixTo_234_dout;
  wire       [15:0]   fixTo_235_dout;
  wire       [15:0]   fixTo_236_dout;
  wire       [15:0]   fixTo_237_dout;
  wire       [15:0]   fixTo_238_dout;
  wire       [15:0]   fixTo_239_dout;
  wire       [15:0]   fixTo_240_dout;
  wire       [15:0]   fixTo_241_dout;
  wire       [15:0]   fixTo_242_dout;
  wire       [15:0]   fixTo_243_dout;
  wire       [15:0]   fixTo_244_dout;
  wire       [15:0]   fixTo_245_dout;
  wire       [15:0]   fixTo_246_dout;
  wire       [15:0]   fixTo_247_dout;
  wire       [15:0]   fixTo_248_dout;
  wire       [15:0]   fixTo_249_dout;
  wire       [15:0]   fixTo_250_dout;
  wire       [15:0]   fixTo_251_dout;
  wire       [15:0]   fixTo_252_dout;
  wire       [15:0]   fixTo_253_dout;
  wire       [15:0]   fixTo_254_dout;
  wire       [15:0]   fixTo_255_dout;
  wire       [15:0]   fixTo_256_dout;
  wire       [15:0]   fixTo_257_dout;
  wire       [15:0]   fixTo_258_dout;
  wire       [15:0]   fixTo_259_dout;
  wire       [15:0]   fixTo_260_dout;
  wire       [15:0]   fixTo_261_dout;
  wire       [15:0]   fixTo_262_dout;
  wire       [15:0]   fixTo_263_dout;
  wire       [15:0]   fixTo_264_dout;
  wire       [15:0]   fixTo_265_dout;
  wire       [15:0]   fixTo_266_dout;
  wire       [15:0]   fixTo_267_dout;
  wire       [15:0]   fixTo_268_dout;
  wire       [15:0]   fixTo_269_dout;
  wire       [15:0]   fixTo_270_dout;
  wire       [15:0]   fixTo_271_dout;
  wire       [15:0]   fixTo_272_dout;
  wire       [15:0]   fixTo_273_dout;
  wire       [15:0]   fixTo_274_dout;
  wire       [15:0]   fixTo_275_dout;
  wire       [15:0]   fixTo_276_dout;
  wire       [15:0]   fixTo_277_dout;
  wire       [15:0]   fixTo_278_dout;
  wire       [15:0]   fixTo_279_dout;
  wire       [15:0]   fixTo_280_dout;
  wire       [15:0]   fixTo_281_dout;
  wire       [15:0]   fixTo_282_dout;
  wire       [15:0]   fixTo_283_dout;
  wire       [15:0]   fixTo_284_dout;
  wire       [15:0]   fixTo_285_dout;
  wire       [15:0]   fixTo_286_dout;
  wire       [15:0]   fixTo_287_dout;
  wire       [15:0]   fixTo_288_dout;
  wire       [15:0]   fixTo_289_dout;
  wire       [15:0]   fixTo_290_dout;
  wire       [15:0]   fixTo_291_dout;
  wire       [15:0]   fixTo_292_dout;
  wire       [15:0]   fixTo_293_dout;
  wire       [15:0]   fixTo_294_dout;
  wire       [15:0]   fixTo_295_dout;
  wire       [15:0]   fixTo_296_dout;
  wire       [15:0]   fixTo_297_dout;
  wire       [15:0]   fixTo_298_dout;
  wire       [15:0]   fixTo_299_dout;
  wire       [15:0]   fixTo_300_dout;
  wire       [15:0]   fixTo_301_dout;
  wire       [15:0]   fixTo_302_dout;
  wire       [15:0]   fixTo_303_dout;
  wire       [15:0]   fixTo_304_dout;
  wire       [15:0]   fixTo_305_dout;
  wire       [15:0]   fixTo_306_dout;
  wire       [15:0]   fixTo_307_dout;
  wire       [15:0]   fixTo_308_dout;
  wire       [15:0]   fixTo_309_dout;
  wire       [15:0]   fixTo_310_dout;
  wire       [15:0]   fixTo_311_dout;
  wire       [15:0]   fixTo_312_dout;
  wire       [15:0]   fixTo_313_dout;
  wire       [15:0]   fixTo_314_dout;
  wire       [15:0]   fixTo_315_dout;
  wire       [15:0]   fixTo_316_dout;
  wire       [15:0]   fixTo_317_dout;
  wire       [15:0]   fixTo_318_dout;
  wire       [15:0]   fixTo_319_dout;
  wire       [15:0]   fixTo_320_dout;
  wire       [15:0]   fixTo_321_dout;
  wire       [15:0]   fixTo_322_dout;
  wire       [15:0]   fixTo_323_dout;
  wire       [15:0]   fixTo_324_dout;
  wire       [15:0]   fixTo_325_dout;
  wire       [15:0]   fixTo_326_dout;
  wire       [15:0]   fixTo_327_dout;
  wire       [15:0]   fixTo_328_dout;
  wire       [15:0]   fixTo_329_dout;
  wire       [15:0]   fixTo_330_dout;
  wire       [15:0]   fixTo_331_dout;
  wire       [15:0]   fixTo_332_dout;
  wire       [15:0]   fixTo_333_dout;
  wire       [15:0]   fixTo_334_dout;
  wire       [15:0]   fixTo_335_dout;
  wire       [15:0]   fixTo_336_dout;
  wire       [15:0]   fixTo_337_dout;
  wire       [15:0]   fixTo_338_dout;
  wire       [15:0]   fixTo_339_dout;
  wire       [15:0]   fixTo_340_dout;
  wire       [15:0]   fixTo_341_dout;
  wire       [15:0]   fixTo_342_dout;
  wire       [15:0]   fixTo_343_dout;
  wire       [15:0]   fixTo_344_dout;
  wire       [15:0]   fixTo_345_dout;
  wire       [15:0]   fixTo_346_dout;
  wire       [15:0]   fixTo_347_dout;
  wire       [15:0]   fixTo_348_dout;
  wire       [15:0]   fixTo_349_dout;
  wire       [15:0]   fixTo_350_dout;
  wire       [15:0]   fixTo_351_dout;
  wire       [15:0]   fixTo_352_dout;
  wire       [15:0]   fixTo_353_dout;
  wire       [15:0]   fixTo_354_dout;
  wire       [15:0]   fixTo_355_dout;
  wire       [15:0]   fixTo_356_dout;
  wire       [15:0]   fixTo_357_dout;
  wire       [15:0]   fixTo_358_dout;
  wire       [15:0]   fixTo_359_dout;
  wire       [15:0]   fixTo_360_dout;
  wire       [15:0]   fixTo_361_dout;
  wire       [15:0]   fixTo_362_dout;
  wire       [15:0]   fixTo_363_dout;
  wire       [15:0]   fixTo_364_dout;
  wire       [15:0]   fixTo_365_dout;
  wire       [15:0]   fixTo_366_dout;
  wire       [15:0]   fixTo_367_dout;
  wire       [15:0]   fixTo_368_dout;
  wire       [15:0]   fixTo_369_dout;
  wire       [15:0]   fixTo_370_dout;
  wire       [15:0]   fixTo_371_dout;
  wire       [15:0]   fixTo_372_dout;
  wire       [15:0]   fixTo_373_dout;
  wire       [15:0]   fixTo_374_dout;
  wire       [15:0]   fixTo_375_dout;
  wire       [15:0]   fixTo_376_dout;
  wire       [15:0]   fixTo_377_dout;
  wire       [15:0]   fixTo_378_dout;
  wire       [15:0]   fixTo_379_dout;
  wire       [15:0]   fixTo_380_dout;
  wire       [15:0]   fixTo_381_dout;
  wire       [15:0]   fixTo_382_dout;
  wire       [15:0]   fixTo_383_dout;
  wire       [15:0]   fixTo_384_dout;
  wire       [15:0]   fixTo_385_dout;
  wire       [15:0]   fixTo_386_dout;
  wire       [15:0]   fixTo_387_dout;
  wire       [15:0]   fixTo_388_dout;
  wire       [15:0]   fixTo_389_dout;
  wire       [15:0]   fixTo_390_dout;
  wire       [15:0]   fixTo_391_dout;
  wire       [15:0]   fixTo_392_dout;
  wire       [15:0]   fixTo_393_dout;
  wire       [15:0]   fixTo_394_dout;
  wire       [15:0]   fixTo_395_dout;
  wire       [15:0]   fixTo_396_dout;
  wire       [15:0]   fixTo_397_dout;
  wire       [15:0]   fixTo_398_dout;
  wire       [15:0]   fixTo_399_dout;
  wire       [15:0]   fixTo_400_dout;
  wire       [15:0]   fixTo_401_dout;
  wire       [15:0]   fixTo_402_dout;
  wire       [15:0]   fixTo_403_dout;
  wire       [15:0]   fixTo_404_dout;
  wire       [15:0]   fixTo_405_dout;
  wire       [15:0]   fixTo_406_dout;
  wire       [15:0]   fixTo_407_dout;
  wire       [15:0]   fixTo_408_dout;
  wire       [15:0]   fixTo_409_dout;
  wire       [15:0]   fixTo_410_dout;
  wire       [15:0]   fixTo_411_dout;
  wire       [15:0]   fixTo_412_dout;
  wire       [15:0]   fixTo_413_dout;
  wire       [15:0]   fixTo_414_dout;
  wire       [15:0]   fixTo_415_dout;
  wire       [15:0]   fixTo_416_dout;
  wire       [15:0]   fixTo_417_dout;
  wire       [15:0]   fixTo_418_dout;
  wire       [15:0]   fixTo_419_dout;
  wire       [15:0]   fixTo_420_dout;
  wire       [15:0]   fixTo_421_dout;
  wire       [15:0]   fixTo_422_dout;
  wire       [15:0]   fixTo_423_dout;
  wire       [15:0]   fixTo_424_dout;
  wire       [15:0]   fixTo_425_dout;
  wire       [15:0]   fixTo_426_dout;
  wire       [15:0]   fixTo_427_dout;
  wire       [15:0]   fixTo_428_dout;
  wire       [15:0]   fixTo_429_dout;
  wire       [15:0]   fixTo_430_dout;
  wire       [15:0]   fixTo_431_dout;
  wire       [15:0]   fixTo_432_dout;
  wire       [15:0]   fixTo_433_dout;
  wire       [15:0]   fixTo_434_dout;
  wire       [15:0]   fixTo_435_dout;
  wire       [15:0]   fixTo_436_dout;
  wire       [15:0]   fixTo_437_dout;
  wire       [15:0]   fixTo_438_dout;
  wire       [15:0]   fixTo_439_dout;
  wire       [15:0]   fixTo_440_dout;
  wire       [15:0]   fixTo_441_dout;
  wire       [15:0]   fixTo_442_dout;
  wire       [15:0]   fixTo_443_dout;
  wire       [15:0]   fixTo_444_dout;
  wire       [15:0]   fixTo_445_dout;
  wire       [15:0]   fixTo_446_dout;
  wire       [15:0]   fixTo_447_dout;
  wire       [15:0]   fixTo_448_dout;
  wire       [15:0]   fixTo_449_dout;
  wire       [15:0]   fixTo_450_dout;
  wire       [15:0]   fixTo_451_dout;
  wire       [15:0]   fixTo_452_dout;
  wire       [15:0]   fixTo_453_dout;
  wire       [15:0]   fixTo_454_dout;
  wire       [15:0]   fixTo_455_dout;
  wire       [15:0]   fixTo_456_dout;
  wire       [15:0]   fixTo_457_dout;
  wire       [15:0]   fixTo_458_dout;
  wire       [15:0]   fixTo_459_dout;
  wire       [15:0]   fixTo_460_dout;
  wire       [15:0]   fixTo_461_dout;
  wire       [15:0]   fixTo_462_dout;
  wire       [15:0]   fixTo_463_dout;
  wire       [15:0]   fixTo_464_dout;
  wire       [15:0]   fixTo_465_dout;
  wire       [15:0]   fixTo_466_dout;
  wire       [15:0]   fixTo_467_dout;
  wire       [15:0]   fixTo_468_dout;
  wire       [15:0]   fixTo_469_dout;
  wire       [15:0]   fixTo_470_dout;
  wire       [15:0]   fixTo_471_dout;
  wire       [15:0]   fixTo_472_dout;
  wire       [15:0]   fixTo_473_dout;
  wire       [15:0]   fixTo_474_dout;
  wire       [15:0]   fixTo_475_dout;
  wire       [15:0]   fixTo_476_dout;
  wire       [15:0]   fixTo_477_dout;
  wire       [15:0]   fixTo_478_dout;
  wire       [15:0]   fixTo_479_dout;
  wire       [15:0]   fixTo_480_dout;
  wire       [15:0]   fixTo_481_dout;
  wire       [15:0]   fixTo_482_dout;
  wire       [15:0]   fixTo_483_dout;
  wire       [15:0]   fixTo_484_dout;
  wire       [15:0]   fixTo_485_dout;
  wire       [15:0]   fixTo_486_dout;
  wire       [15:0]   fixTo_487_dout;
  wire       [15:0]   fixTo_488_dout;
  wire       [15:0]   fixTo_489_dout;
  wire       [15:0]   fixTo_490_dout;
  wire       [15:0]   fixTo_491_dout;
  wire       [15:0]   fixTo_492_dout;
  wire       [15:0]   fixTo_493_dout;
  wire       [15:0]   fixTo_494_dout;
  wire       [15:0]   fixTo_495_dout;
  wire       [15:0]   fixTo_496_dout;
  wire       [15:0]   fixTo_497_dout;
  wire       [15:0]   fixTo_498_dout;
  wire       [15:0]   fixTo_499_dout;
  wire       [15:0]   fixTo_500_dout;
  wire       [15:0]   fixTo_501_dout;
  wire       [15:0]   fixTo_502_dout;
  wire       [15:0]   fixTo_503_dout;
  wire       [15:0]   fixTo_504_dout;
  wire       [15:0]   fixTo_505_dout;
  wire       [15:0]   fixTo_506_dout;
  wire       [15:0]   fixTo_507_dout;
  wire       [15:0]   fixTo_508_dout;
  wire       [15:0]   fixTo_509_dout;
  wire       [15:0]   fixTo_510_dout;
  wire       [15:0]   fixTo_511_dout;
  wire       [15:0]   fixTo_512_dout;
  wire       [15:0]   fixTo_513_dout;
  wire       [15:0]   fixTo_514_dout;
  wire       [15:0]   fixTo_515_dout;
  wire       [15:0]   fixTo_516_dout;
  wire       [15:0]   fixTo_517_dout;
  wire       [15:0]   fixTo_518_dout;
  wire       [15:0]   fixTo_519_dout;
  wire       [15:0]   fixTo_520_dout;
  wire       [15:0]   fixTo_521_dout;
  wire       [15:0]   fixTo_522_dout;
  wire       [15:0]   fixTo_523_dout;
  wire       [15:0]   fixTo_524_dout;
  wire       [15:0]   fixTo_525_dout;
  wire       [15:0]   fixTo_526_dout;
  wire       [15:0]   fixTo_527_dout;
  wire       [15:0]   fixTo_528_dout;
  wire       [15:0]   fixTo_529_dout;
  wire       [15:0]   fixTo_530_dout;
  wire       [15:0]   fixTo_531_dout;
  wire       [15:0]   fixTo_532_dout;
  wire       [15:0]   fixTo_533_dout;
  wire       [15:0]   fixTo_534_dout;
  wire       [15:0]   fixTo_535_dout;
  wire       [15:0]   fixTo_536_dout;
  wire       [15:0]   fixTo_537_dout;
  wire       [15:0]   fixTo_538_dout;
  wire       [15:0]   fixTo_539_dout;
  wire       [15:0]   fixTo_540_dout;
  wire       [15:0]   fixTo_541_dout;
  wire       [15:0]   fixTo_542_dout;
  wire       [15:0]   fixTo_543_dout;
  wire       [15:0]   fixTo_544_dout;
  wire       [15:0]   fixTo_545_dout;
  wire       [15:0]   fixTo_546_dout;
  wire       [15:0]   fixTo_547_dout;
  wire       [15:0]   fixTo_548_dout;
  wire       [15:0]   fixTo_549_dout;
  wire       [15:0]   fixTo_550_dout;
  wire       [15:0]   fixTo_551_dout;
  wire       [15:0]   fixTo_552_dout;
  wire       [15:0]   fixTo_553_dout;
  wire       [15:0]   fixTo_554_dout;
  wire       [15:0]   fixTo_555_dout;
  wire       [15:0]   fixTo_556_dout;
  wire       [15:0]   fixTo_557_dout;
  wire       [15:0]   fixTo_558_dout;
  wire       [15:0]   fixTo_559_dout;
  wire       [15:0]   fixTo_560_dout;
  wire       [15:0]   fixTo_561_dout;
  wire       [15:0]   fixTo_562_dout;
  wire       [15:0]   fixTo_563_dout;
  wire       [15:0]   fixTo_564_dout;
  wire       [15:0]   fixTo_565_dout;
  wire       [15:0]   fixTo_566_dout;
  wire       [15:0]   fixTo_567_dout;
  wire       [15:0]   fixTo_568_dout;
  wire       [15:0]   fixTo_569_dout;
  wire       [15:0]   fixTo_570_dout;
  wire       [15:0]   fixTo_571_dout;
  wire       [15:0]   fixTo_572_dout;
  wire       [15:0]   fixTo_573_dout;
  wire       [15:0]   fixTo_574_dout;
  wire       [15:0]   fixTo_575_dout;
  wire       [15:0]   fixTo_576_dout;
  wire       [15:0]   fixTo_577_dout;
  wire       [15:0]   fixTo_578_dout;
  wire       [15:0]   fixTo_579_dout;
  wire       [15:0]   fixTo_580_dout;
  wire       [15:0]   fixTo_581_dout;
  wire       [15:0]   fixTo_582_dout;
  wire       [15:0]   fixTo_583_dout;
  wire       [15:0]   fixTo_584_dout;
  wire       [15:0]   fixTo_585_dout;
  wire       [15:0]   fixTo_586_dout;
  wire       [15:0]   fixTo_587_dout;
  wire       [15:0]   fixTo_588_dout;
  wire       [15:0]   fixTo_589_dout;
  wire       [15:0]   fixTo_590_dout;
  wire       [15:0]   fixTo_591_dout;
  wire       [15:0]   fixTo_592_dout;
  wire       [15:0]   fixTo_593_dout;
  wire       [15:0]   fixTo_594_dout;
  wire       [15:0]   fixTo_595_dout;
  wire       [15:0]   fixTo_596_dout;
  wire       [15:0]   fixTo_597_dout;
  wire       [15:0]   fixTo_598_dout;
  wire       [15:0]   fixTo_599_dout;
  wire       [15:0]   fixTo_600_dout;
  wire       [15:0]   fixTo_601_dout;
  wire       [15:0]   fixTo_602_dout;
  wire       [15:0]   fixTo_603_dout;
  wire       [15:0]   fixTo_604_dout;
  wire       [15:0]   fixTo_605_dout;
  wire       [15:0]   fixTo_606_dout;
  wire       [15:0]   fixTo_607_dout;
  wire       [15:0]   fixTo_608_dout;
  wire       [15:0]   fixTo_609_dout;
  wire       [15:0]   fixTo_610_dout;
  wire       [15:0]   fixTo_611_dout;
  wire       [15:0]   fixTo_612_dout;
  wire       [15:0]   fixTo_613_dout;
  wire       [15:0]   fixTo_614_dout;
  wire       [15:0]   fixTo_615_dout;
  wire       [15:0]   fixTo_616_dout;
  wire       [15:0]   fixTo_617_dout;
  wire       [15:0]   fixTo_618_dout;
  wire       [15:0]   fixTo_619_dout;
  wire       [15:0]   fixTo_620_dout;
  wire       [15:0]   fixTo_621_dout;
  wire       [15:0]   fixTo_622_dout;
  wire       [15:0]   fixTo_623_dout;
  wire       [15:0]   fixTo_624_dout;
  wire       [15:0]   fixTo_625_dout;
  wire       [15:0]   fixTo_626_dout;
  wire       [15:0]   fixTo_627_dout;
  wire       [15:0]   fixTo_628_dout;
  wire       [15:0]   fixTo_629_dout;
  wire       [15:0]   fixTo_630_dout;
  wire       [15:0]   fixTo_631_dout;
  wire       [15:0]   fixTo_632_dout;
  wire       [15:0]   fixTo_633_dout;
  wire       [15:0]   fixTo_634_dout;
  wire       [15:0]   fixTo_635_dout;
  wire       [15:0]   fixTo_636_dout;
  wire       [15:0]   fixTo_637_dout;
  wire       [15:0]   fixTo_638_dout;
  wire       [15:0]   fixTo_639_dout;
  wire       [15:0]   fixTo_640_dout;
  wire       [15:0]   fixTo_641_dout;
  wire       [15:0]   fixTo_642_dout;
  wire       [15:0]   fixTo_643_dout;
  wire       [15:0]   fixTo_644_dout;
  wire       [15:0]   fixTo_645_dout;
  wire       [15:0]   fixTo_646_dout;
  wire       [15:0]   fixTo_647_dout;
  wire       [15:0]   fixTo_648_dout;
  wire       [15:0]   fixTo_649_dout;
  wire       [15:0]   fixTo_650_dout;
  wire       [15:0]   fixTo_651_dout;
  wire       [15:0]   fixTo_652_dout;
  wire       [15:0]   fixTo_653_dout;
  wire       [15:0]   fixTo_654_dout;
  wire       [15:0]   fixTo_655_dout;
  wire       [15:0]   fixTo_656_dout;
  wire       [15:0]   fixTo_657_dout;
  wire       [15:0]   fixTo_658_dout;
  wire       [15:0]   fixTo_659_dout;
  wire       [15:0]   fixTo_660_dout;
  wire       [15:0]   fixTo_661_dout;
  wire       [15:0]   fixTo_662_dout;
  wire       [15:0]   fixTo_663_dout;
  wire       [15:0]   fixTo_664_dout;
  wire       [15:0]   fixTo_665_dout;
  wire       [15:0]   fixTo_666_dout;
  wire       [15:0]   fixTo_667_dout;
  wire       [15:0]   fixTo_668_dout;
  wire       [15:0]   fixTo_669_dout;
  wire       [15:0]   fixTo_670_dout;
  wire       [15:0]   fixTo_671_dout;
  wire       [15:0]   fixTo_672_dout;
  wire       [15:0]   fixTo_673_dout;
  wire       [15:0]   fixTo_674_dout;
  wire       [15:0]   fixTo_675_dout;
  wire       [15:0]   fixTo_676_dout;
  wire       [15:0]   fixTo_677_dout;
  wire       [15:0]   fixTo_678_dout;
  wire       [15:0]   fixTo_679_dout;
  wire       [15:0]   fixTo_680_dout;
  wire       [15:0]   fixTo_681_dout;
  wire       [15:0]   fixTo_682_dout;
  wire       [15:0]   fixTo_683_dout;
  wire       [15:0]   fixTo_684_dout;
  wire       [15:0]   fixTo_685_dout;
  wire       [15:0]   fixTo_686_dout;
  wire       [15:0]   fixTo_687_dout;
  wire       [15:0]   fixTo_688_dout;
  wire       [15:0]   fixTo_689_dout;
  wire       [15:0]   fixTo_690_dout;
  wire       [15:0]   fixTo_691_dout;
  wire       [15:0]   fixTo_692_dout;
  wire       [15:0]   fixTo_693_dout;
  wire       [15:0]   fixTo_694_dout;
  wire       [15:0]   fixTo_695_dout;
  wire       [15:0]   fixTo_696_dout;
  wire       [15:0]   fixTo_697_dout;
  wire       [15:0]   fixTo_698_dout;
  wire       [15:0]   fixTo_699_dout;
  wire       [15:0]   fixTo_700_dout;
  wire       [15:0]   fixTo_701_dout;
  wire       [15:0]   fixTo_702_dout;
  wire       [15:0]   fixTo_703_dout;
  wire       [15:0]   fixTo_704_dout;
  wire       [15:0]   fixTo_705_dout;
  wire       [15:0]   fixTo_706_dout;
  wire       [15:0]   fixTo_707_dout;
  wire       [15:0]   fixTo_708_dout;
  wire       [15:0]   fixTo_709_dout;
  wire       [15:0]   fixTo_710_dout;
  wire       [15:0]   fixTo_711_dout;
  wire       [15:0]   fixTo_712_dout;
  wire       [15:0]   fixTo_713_dout;
  wire       [15:0]   fixTo_714_dout;
  wire       [15:0]   fixTo_715_dout;
  wire       [15:0]   fixTo_716_dout;
  wire       [15:0]   fixTo_717_dout;
  wire       [15:0]   fixTo_718_dout;
  wire       [15:0]   fixTo_719_dout;
  wire       [15:0]   fixTo_720_dout;
  wire       [15:0]   fixTo_721_dout;
  wire       [15:0]   fixTo_722_dout;
  wire       [15:0]   fixTo_723_dout;
  wire       [15:0]   fixTo_724_dout;
  wire       [15:0]   fixTo_725_dout;
  wire       [15:0]   fixTo_726_dout;
  wire       [15:0]   fixTo_727_dout;
  wire       [15:0]   fixTo_728_dout;
  wire       [15:0]   fixTo_729_dout;
  wire       [15:0]   fixTo_730_dout;
  wire       [15:0]   fixTo_731_dout;
  wire       [15:0]   fixTo_732_dout;
  wire       [15:0]   fixTo_733_dout;
  wire       [15:0]   fixTo_734_dout;
  wire       [15:0]   fixTo_735_dout;
  wire       [15:0]   fixTo_736_dout;
  wire       [15:0]   fixTo_737_dout;
  wire       [15:0]   fixTo_738_dout;
  wire       [15:0]   fixTo_739_dout;
  wire       [15:0]   fixTo_740_dout;
  wire       [15:0]   fixTo_741_dout;
  wire       [15:0]   fixTo_742_dout;
  wire       [15:0]   fixTo_743_dout;
  wire       [15:0]   fixTo_744_dout;
  wire       [15:0]   fixTo_745_dout;
  wire       [15:0]   fixTo_746_dout;
  wire       [15:0]   fixTo_747_dout;
  wire       [15:0]   fixTo_748_dout;
  wire       [15:0]   fixTo_749_dout;
  wire       [15:0]   fixTo_750_dout;
  wire       [15:0]   fixTo_751_dout;
  wire       [15:0]   fixTo_752_dout;
  wire       [15:0]   fixTo_753_dout;
  wire       [15:0]   fixTo_754_dout;
  wire       [15:0]   fixTo_755_dout;
  wire       [15:0]   fixTo_756_dout;
  wire       [15:0]   fixTo_757_dout;
  wire       [15:0]   fixTo_758_dout;
  wire       [15:0]   fixTo_759_dout;
  wire       [15:0]   fixTo_760_dout;
  wire       [15:0]   fixTo_761_dout;
  wire       [15:0]   fixTo_762_dout;
  wire       [15:0]   fixTo_763_dout;
  wire       [15:0]   fixTo_764_dout;
  wire       [15:0]   fixTo_765_dout;
  wire       [15:0]   fixTo_766_dout;
  wire       [15:0]   fixTo_767_dout;
  wire       [15:0]   fixTo_768_dout;
  wire       [15:0]   fixTo_769_dout;
  wire       [15:0]   fixTo_770_dout;
  wire       [15:0]   fixTo_771_dout;
  wire       [15:0]   fixTo_772_dout;
  wire       [15:0]   fixTo_773_dout;
  wire       [15:0]   fixTo_774_dout;
  wire       [15:0]   fixTo_775_dout;
  wire       [15:0]   fixTo_776_dout;
  wire       [15:0]   fixTo_777_dout;
  wire       [15:0]   fixTo_778_dout;
  wire       [15:0]   fixTo_779_dout;
  wire       [15:0]   fixTo_780_dout;
  wire       [15:0]   fixTo_781_dout;
  wire       [15:0]   fixTo_782_dout;
  wire       [15:0]   fixTo_783_dout;
  wire       [15:0]   fixTo_784_dout;
  wire       [15:0]   fixTo_785_dout;
  wire       [15:0]   fixTo_786_dout;
  wire       [15:0]   fixTo_787_dout;
  wire       [15:0]   fixTo_788_dout;
  wire       [15:0]   fixTo_789_dout;
  wire       [15:0]   fixTo_790_dout;
  wire       [15:0]   fixTo_791_dout;
  wire       [15:0]   fixTo_792_dout;
  wire       [15:0]   fixTo_793_dout;
  wire       [15:0]   fixTo_794_dout;
  wire       [15:0]   fixTo_795_dout;
  wire       [15:0]   fixTo_796_dout;
  wire       [15:0]   fixTo_797_dout;
  wire       [15:0]   fixTo_798_dout;
  wire       [15:0]   fixTo_799_dout;
  wire       [15:0]   fixTo_800_dout;
  wire       [15:0]   fixTo_801_dout;
  wire       [15:0]   fixTo_802_dout;
  wire       [15:0]   fixTo_803_dout;
  wire       [15:0]   fixTo_804_dout;
  wire       [15:0]   fixTo_805_dout;
  wire       [15:0]   fixTo_806_dout;
  wire       [15:0]   fixTo_807_dout;
  wire       [15:0]   fixTo_808_dout;
  wire       [15:0]   fixTo_809_dout;
  wire       [15:0]   fixTo_810_dout;
  wire       [15:0]   fixTo_811_dout;
  wire       [15:0]   fixTo_812_dout;
  wire       [15:0]   fixTo_813_dout;
  wire       [15:0]   fixTo_814_dout;
  wire       [15:0]   fixTo_815_dout;
  wire       [15:0]   fixTo_816_dout;
  wire       [15:0]   fixTo_817_dout;
  wire       [15:0]   fixTo_818_dout;
  wire       [15:0]   fixTo_819_dout;
  wire       [15:0]   fixTo_820_dout;
  wire       [15:0]   fixTo_821_dout;
  wire       [15:0]   fixTo_822_dout;
  wire       [15:0]   fixTo_823_dout;
  wire       [15:0]   fixTo_824_dout;
  wire       [15:0]   fixTo_825_dout;
  wire       [15:0]   fixTo_826_dout;
  wire       [15:0]   fixTo_827_dout;
  wire       [15:0]   fixTo_828_dout;
  wire       [15:0]   fixTo_829_dout;
  wire       [15:0]   fixTo_830_dout;
  wire       [15:0]   fixTo_831_dout;
  wire       [15:0]   fixTo_832_dout;
  wire       [15:0]   fixTo_833_dout;
  wire       [15:0]   fixTo_834_dout;
  wire       [15:0]   fixTo_835_dout;
  wire       [15:0]   fixTo_836_dout;
  wire       [15:0]   fixTo_837_dout;
  wire       [15:0]   fixTo_838_dout;
  wire       [15:0]   fixTo_839_dout;
  wire       [15:0]   fixTo_840_dout;
  wire       [15:0]   fixTo_841_dout;
  wire       [15:0]   fixTo_842_dout;
  wire       [15:0]   fixTo_843_dout;
  wire       [15:0]   fixTo_844_dout;
  wire       [15:0]   fixTo_845_dout;
  wire       [15:0]   fixTo_846_dout;
  wire       [15:0]   fixTo_847_dout;
  wire       [15:0]   fixTo_848_dout;
  wire       [15:0]   fixTo_849_dout;
  wire       [15:0]   fixTo_850_dout;
  wire       [15:0]   fixTo_851_dout;
  wire       [15:0]   fixTo_852_dout;
  wire       [15:0]   fixTo_853_dout;
  wire       [15:0]   fixTo_854_dout;
  wire       [15:0]   fixTo_855_dout;
  wire       [15:0]   fixTo_856_dout;
  wire       [15:0]   fixTo_857_dout;
  wire       [15:0]   fixTo_858_dout;
  wire       [15:0]   fixTo_859_dout;
  wire       [15:0]   fixTo_860_dout;
  wire       [15:0]   fixTo_861_dout;
  wire       [15:0]   fixTo_862_dout;
  wire       [15:0]   fixTo_863_dout;
  wire       [15:0]   fixTo_864_dout;
  wire       [15:0]   fixTo_865_dout;
  wire       [15:0]   fixTo_866_dout;
  wire       [15:0]   fixTo_867_dout;
  wire       [15:0]   fixTo_868_dout;
  wire       [15:0]   fixTo_869_dout;
  wire       [15:0]   fixTo_870_dout;
  wire       [15:0]   fixTo_871_dout;
  wire       [15:0]   fixTo_872_dout;
  wire       [15:0]   fixTo_873_dout;
  wire       [15:0]   fixTo_874_dout;
  wire       [15:0]   fixTo_875_dout;
  wire       [15:0]   fixTo_876_dout;
  wire       [15:0]   fixTo_877_dout;
  wire       [15:0]   fixTo_878_dout;
  wire       [15:0]   fixTo_879_dout;
  wire       [15:0]   fixTo_880_dout;
  wire       [15:0]   fixTo_881_dout;
  wire       [15:0]   fixTo_882_dout;
  wire       [15:0]   fixTo_883_dout;
  wire       [15:0]   fixTo_884_dout;
  wire       [15:0]   fixTo_885_dout;
  wire       [15:0]   fixTo_886_dout;
  wire       [15:0]   fixTo_887_dout;
  wire       [15:0]   fixTo_888_dout;
  wire       [15:0]   fixTo_889_dout;
  wire       [15:0]   fixTo_890_dout;
  wire       [15:0]   fixTo_891_dout;
  wire       [15:0]   fixTo_892_dout;
  wire       [15:0]   fixTo_893_dout;
  wire       [15:0]   fixTo_894_dout;
  wire       [15:0]   fixTo_895_dout;
  wire       [0:0]    _zz_2689;
  wire       [2:0]    _zz_2690;
  wire       [31:0]   _zz_2691;
  wire       [31:0]   _zz_2692;
  wire       [15:0]   _zz_2693;
  wire       [31:0]   _zz_2694;
  wire       [31:0]   _zz_2695;
  wire       [15:0]   _zz_2696;
  wire       [15:0]   _zz_2697;
  wire       [15:0]   _zz_2698;
  wire       [15:0]   _zz_2699;
  wire       [15:0]   _zz_2700;
  wire       [15:0]   _zz_2701;
  wire       [15:0]   _zz_2702;
  wire       [15:0]   _zz_2703;
  wire       [15:0]   _zz_2704;
  wire       [15:0]   _zz_2705;
  wire       [15:0]   _zz_2706;
  wire       [15:0]   _zz_2707;
  wire       [15:0]   _zz_2708;
  wire       [15:0]   _zz_2709;
  wire       [15:0]   _zz_2710;
  wire       [15:0]   _zz_2711;
  wire       [15:0]   _zz_2712;
  wire       [31:0]   _zz_2713;
  wire       [31:0]   _zz_2714;
  wire       [15:0]   _zz_2715;
  wire       [31:0]   _zz_2716;
  wire       [31:0]   _zz_2717;
  wire       [15:0]   _zz_2718;
  wire       [15:0]   _zz_2719;
  wire       [15:0]   _zz_2720;
  wire       [15:0]   _zz_2721;
  wire       [15:0]   _zz_2722;
  wire       [15:0]   _zz_2723;
  wire       [15:0]   _zz_2724;
  wire       [15:0]   _zz_2725;
  wire       [15:0]   _zz_2726;
  wire       [15:0]   _zz_2727;
  wire       [15:0]   _zz_2728;
  wire       [15:0]   _zz_2729;
  wire       [15:0]   _zz_2730;
  wire       [15:0]   _zz_2731;
  wire       [15:0]   _zz_2732;
  wire       [15:0]   _zz_2733;
  wire       [15:0]   _zz_2734;
  wire       [31:0]   _zz_2735;
  wire       [31:0]   _zz_2736;
  wire       [15:0]   _zz_2737;
  wire       [31:0]   _zz_2738;
  wire       [31:0]   _zz_2739;
  wire       [15:0]   _zz_2740;
  wire       [15:0]   _zz_2741;
  wire       [15:0]   _zz_2742;
  wire       [15:0]   _zz_2743;
  wire       [15:0]   _zz_2744;
  wire       [15:0]   _zz_2745;
  wire       [15:0]   _zz_2746;
  wire       [15:0]   _zz_2747;
  wire       [15:0]   _zz_2748;
  wire       [15:0]   _zz_2749;
  wire       [15:0]   _zz_2750;
  wire       [15:0]   _zz_2751;
  wire       [15:0]   _zz_2752;
  wire       [15:0]   _zz_2753;
  wire       [15:0]   _zz_2754;
  wire       [15:0]   _zz_2755;
  wire       [15:0]   _zz_2756;
  wire       [31:0]   _zz_2757;
  wire       [31:0]   _zz_2758;
  wire       [15:0]   _zz_2759;
  wire       [31:0]   _zz_2760;
  wire       [31:0]   _zz_2761;
  wire       [15:0]   _zz_2762;
  wire       [15:0]   _zz_2763;
  wire       [15:0]   _zz_2764;
  wire       [15:0]   _zz_2765;
  wire       [15:0]   _zz_2766;
  wire       [15:0]   _zz_2767;
  wire       [15:0]   _zz_2768;
  wire       [15:0]   _zz_2769;
  wire       [15:0]   _zz_2770;
  wire       [15:0]   _zz_2771;
  wire       [15:0]   _zz_2772;
  wire       [15:0]   _zz_2773;
  wire       [15:0]   _zz_2774;
  wire       [15:0]   _zz_2775;
  wire       [15:0]   _zz_2776;
  wire       [15:0]   _zz_2777;
  wire       [15:0]   _zz_2778;
  wire       [31:0]   _zz_2779;
  wire       [31:0]   _zz_2780;
  wire       [15:0]   _zz_2781;
  wire       [31:0]   _zz_2782;
  wire       [31:0]   _zz_2783;
  wire       [15:0]   _zz_2784;
  wire       [15:0]   _zz_2785;
  wire       [15:0]   _zz_2786;
  wire       [15:0]   _zz_2787;
  wire       [15:0]   _zz_2788;
  wire       [15:0]   _zz_2789;
  wire       [15:0]   _zz_2790;
  wire       [15:0]   _zz_2791;
  wire       [15:0]   _zz_2792;
  wire       [15:0]   _zz_2793;
  wire       [15:0]   _zz_2794;
  wire       [15:0]   _zz_2795;
  wire       [15:0]   _zz_2796;
  wire       [15:0]   _zz_2797;
  wire       [15:0]   _zz_2798;
  wire       [15:0]   _zz_2799;
  wire       [15:0]   _zz_2800;
  wire       [31:0]   _zz_2801;
  wire       [31:0]   _zz_2802;
  wire       [15:0]   _zz_2803;
  wire       [31:0]   _zz_2804;
  wire       [31:0]   _zz_2805;
  wire       [15:0]   _zz_2806;
  wire       [15:0]   _zz_2807;
  wire       [15:0]   _zz_2808;
  wire       [15:0]   _zz_2809;
  wire       [15:0]   _zz_2810;
  wire       [15:0]   _zz_2811;
  wire       [15:0]   _zz_2812;
  wire       [15:0]   _zz_2813;
  wire       [15:0]   _zz_2814;
  wire       [15:0]   _zz_2815;
  wire       [15:0]   _zz_2816;
  wire       [15:0]   _zz_2817;
  wire       [15:0]   _zz_2818;
  wire       [15:0]   _zz_2819;
  wire       [15:0]   _zz_2820;
  wire       [15:0]   _zz_2821;
  wire       [15:0]   _zz_2822;
  wire       [31:0]   _zz_2823;
  wire       [31:0]   _zz_2824;
  wire       [15:0]   _zz_2825;
  wire       [31:0]   _zz_2826;
  wire       [31:0]   _zz_2827;
  wire       [15:0]   _zz_2828;
  wire       [15:0]   _zz_2829;
  wire       [15:0]   _zz_2830;
  wire       [15:0]   _zz_2831;
  wire       [15:0]   _zz_2832;
  wire       [15:0]   _zz_2833;
  wire       [15:0]   _zz_2834;
  wire       [15:0]   _zz_2835;
  wire       [15:0]   _zz_2836;
  wire       [15:0]   _zz_2837;
  wire       [15:0]   _zz_2838;
  wire       [15:0]   _zz_2839;
  wire       [15:0]   _zz_2840;
  wire       [15:0]   _zz_2841;
  wire       [15:0]   _zz_2842;
  wire       [15:0]   _zz_2843;
  wire       [15:0]   _zz_2844;
  wire       [31:0]   _zz_2845;
  wire       [31:0]   _zz_2846;
  wire       [15:0]   _zz_2847;
  wire       [31:0]   _zz_2848;
  wire       [31:0]   _zz_2849;
  wire       [15:0]   _zz_2850;
  wire       [15:0]   _zz_2851;
  wire       [15:0]   _zz_2852;
  wire       [15:0]   _zz_2853;
  wire       [15:0]   _zz_2854;
  wire       [15:0]   _zz_2855;
  wire       [15:0]   _zz_2856;
  wire       [15:0]   _zz_2857;
  wire       [15:0]   _zz_2858;
  wire       [15:0]   _zz_2859;
  wire       [15:0]   _zz_2860;
  wire       [15:0]   _zz_2861;
  wire       [15:0]   _zz_2862;
  wire       [15:0]   _zz_2863;
  wire       [15:0]   _zz_2864;
  wire       [15:0]   _zz_2865;
  wire       [15:0]   _zz_2866;
  wire       [31:0]   _zz_2867;
  wire       [31:0]   _zz_2868;
  wire       [15:0]   _zz_2869;
  wire       [31:0]   _zz_2870;
  wire       [31:0]   _zz_2871;
  wire       [15:0]   _zz_2872;
  wire       [15:0]   _zz_2873;
  wire       [15:0]   _zz_2874;
  wire       [15:0]   _zz_2875;
  wire       [15:0]   _zz_2876;
  wire       [15:0]   _zz_2877;
  wire       [15:0]   _zz_2878;
  wire       [15:0]   _zz_2879;
  wire       [15:0]   _zz_2880;
  wire       [15:0]   _zz_2881;
  wire       [15:0]   _zz_2882;
  wire       [15:0]   _zz_2883;
  wire       [15:0]   _zz_2884;
  wire       [15:0]   _zz_2885;
  wire       [15:0]   _zz_2886;
  wire       [15:0]   _zz_2887;
  wire       [15:0]   _zz_2888;
  wire       [31:0]   _zz_2889;
  wire       [31:0]   _zz_2890;
  wire       [15:0]   _zz_2891;
  wire       [31:0]   _zz_2892;
  wire       [31:0]   _zz_2893;
  wire       [15:0]   _zz_2894;
  wire       [15:0]   _zz_2895;
  wire       [15:0]   _zz_2896;
  wire       [15:0]   _zz_2897;
  wire       [15:0]   _zz_2898;
  wire       [15:0]   _zz_2899;
  wire       [15:0]   _zz_2900;
  wire       [15:0]   _zz_2901;
  wire       [15:0]   _zz_2902;
  wire       [15:0]   _zz_2903;
  wire       [15:0]   _zz_2904;
  wire       [15:0]   _zz_2905;
  wire       [15:0]   _zz_2906;
  wire       [15:0]   _zz_2907;
  wire       [15:0]   _zz_2908;
  wire       [15:0]   _zz_2909;
  wire       [15:0]   _zz_2910;
  wire       [31:0]   _zz_2911;
  wire       [31:0]   _zz_2912;
  wire       [15:0]   _zz_2913;
  wire       [31:0]   _zz_2914;
  wire       [31:0]   _zz_2915;
  wire       [15:0]   _zz_2916;
  wire       [15:0]   _zz_2917;
  wire       [15:0]   _zz_2918;
  wire       [15:0]   _zz_2919;
  wire       [15:0]   _zz_2920;
  wire       [15:0]   _zz_2921;
  wire       [15:0]   _zz_2922;
  wire       [15:0]   _zz_2923;
  wire       [15:0]   _zz_2924;
  wire       [15:0]   _zz_2925;
  wire       [15:0]   _zz_2926;
  wire       [15:0]   _zz_2927;
  wire       [15:0]   _zz_2928;
  wire       [15:0]   _zz_2929;
  wire       [15:0]   _zz_2930;
  wire       [15:0]   _zz_2931;
  wire       [15:0]   _zz_2932;
  wire       [31:0]   _zz_2933;
  wire       [31:0]   _zz_2934;
  wire       [15:0]   _zz_2935;
  wire       [31:0]   _zz_2936;
  wire       [31:0]   _zz_2937;
  wire       [15:0]   _zz_2938;
  wire       [15:0]   _zz_2939;
  wire       [15:0]   _zz_2940;
  wire       [15:0]   _zz_2941;
  wire       [15:0]   _zz_2942;
  wire       [15:0]   _zz_2943;
  wire       [15:0]   _zz_2944;
  wire       [15:0]   _zz_2945;
  wire       [15:0]   _zz_2946;
  wire       [15:0]   _zz_2947;
  wire       [15:0]   _zz_2948;
  wire       [15:0]   _zz_2949;
  wire       [15:0]   _zz_2950;
  wire       [15:0]   _zz_2951;
  wire       [15:0]   _zz_2952;
  wire       [15:0]   _zz_2953;
  wire       [15:0]   _zz_2954;
  wire       [31:0]   _zz_2955;
  wire       [31:0]   _zz_2956;
  wire       [15:0]   _zz_2957;
  wire       [31:0]   _zz_2958;
  wire       [31:0]   _zz_2959;
  wire       [15:0]   _zz_2960;
  wire       [15:0]   _zz_2961;
  wire       [15:0]   _zz_2962;
  wire       [15:0]   _zz_2963;
  wire       [15:0]   _zz_2964;
  wire       [15:0]   _zz_2965;
  wire       [15:0]   _zz_2966;
  wire       [15:0]   _zz_2967;
  wire       [15:0]   _zz_2968;
  wire       [15:0]   _zz_2969;
  wire       [15:0]   _zz_2970;
  wire       [15:0]   _zz_2971;
  wire       [15:0]   _zz_2972;
  wire       [15:0]   _zz_2973;
  wire       [15:0]   _zz_2974;
  wire       [15:0]   _zz_2975;
  wire       [15:0]   _zz_2976;
  wire       [31:0]   _zz_2977;
  wire       [31:0]   _zz_2978;
  wire       [15:0]   _zz_2979;
  wire       [31:0]   _zz_2980;
  wire       [31:0]   _zz_2981;
  wire       [15:0]   _zz_2982;
  wire       [15:0]   _zz_2983;
  wire       [15:0]   _zz_2984;
  wire       [15:0]   _zz_2985;
  wire       [15:0]   _zz_2986;
  wire       [15:0]   _zz_2987;
  wire       [15:0]   _zz_2988;
  wire       [15:0]   _zz_2989;
  wire       [15:0]   _zz_2990;
  wire       [15:0]   _zz_2991;
  wire       [15:0]   _zz_2992;
  wire       [15:0]   _zz_2993;
  wire       [15:0]   _zz_2994;
  wire       [15:0]   _zz_2995;
  wire       [15:0]   _zz_2996;
  wire       [15:0]   _zz_2997;
  wire       [15:0]   _zz_2998;
  wire       [31:0]   _zz_2999;
  wire       [31:0]   _zz_3000;
  wire       [15:0]   _zz_3001;
  wire       [31:0]   _zz_3002;
  wire       [31:0]   _zz_3003;
  wire       [15:0]   _zz_3004;
  wire       [15:0]   _zz_3005;
  wire       [15:0]   _zz_3006;
  wire       [15:0]   _zz_3007;
  wire       [15:0]   _zz_3008;
  wire       [15:0]   _zz_3009;
  wire       [15:0]   _zz_3010;
  wire       [15:0]   _zz_3011;
  wire       [15:0]   _zz_3012;
  wire       [15:0]   _zz_3013;
  wire       [15:0]   _zz_3014;
  wire       [15:0]   _zz_3015;
  wire       [15:0]   _zz_3016;
  wire       [15:0]   _zz_3017;
  wire       [15:0]   _zz_3018;
  wire       [15:0]   _zz_3019;
  wire       [15:0]   _zz_3020;
  wire       [31:0]   _zz_3021;
  wire       [31:0]   _zz_3022;
  wire       [15:0]   _zz_3023;
  wire       [31:0]   _zz_3024;
  wire       [31:0]   _zz_3025;
  wire       [15:0]   _zz_3026;
  wire       [15:0]   _zz_3027;
  wire       [15:0]   _zz_3028;
  wire       [15:0]   _zz_3029;
  wire       [15:0]   _zz_3030;
  wire       [15:0]   _zz_3031;
  wire       [15:0]   _zz_3032;
  wire       [15:0]   _zz_3033;
  wire       [15:0]   _zz_3034;
  wire       [15:0]   _zz_3035;
  wire       [15:0]   _zz_3036;
  wire       [15:0]   _zz_3037;
  wire       [15:0]   _zz_3038;
  wire       [15:0]   _zz_3039;
  wire       [15:0]   _zz_3040;
  wire       [15:0]   _zz_3041;
  wire       [15:0]   _zz_3042;
  wire       [31:0]   _zz_3043;
  wire       [31:0]   _zz_3044;
  wire       [15:0]   _zz_3045;
  wire       [31:0]   _zz_3046;
  wire       [31:0]   _zz_3047;
  wire       [15:0]   _zz_3048;
  wire       [15:0]   _zz_3049;
  wire       [15:0]   _zz_3050;
  wire       [15:0]   _zz_3051;
  wire       [15:0]   _zz_3052;
  wire       [15:0]   _zz_3053;
  wire       [15:0]   _zz_3054;
  wire       [15:0]   _zz_3055;
  wire       [15:0]   _zz_3056;
  wire       [15:0]   _zz_3057;
  wire       [15:0]   _zz_3058;
  wire       [15:0]   _zz_3059;
  wire       [15:0]   _zz_3060;
  wire       [15:0]   _zz_3061;
  wire       [15:0]   _zz_3062;
  wire       [15:0]   _zz_3063;
  wire       [15:0]   _zz_3064;
  wire       [31:0]   _zz_3065;
  wire       [31:0]   _zz_3066;
  wire       [15:0]   _zz_3067;
  wire       [31:0]   _zz_3068;
  wire       [31:0]   _zz_3069;
  wire       [15:0]   _zz_3070;
  wire       [15:0]   _zz_3071;
  wire       [15:0]   _zz_3072;
  wire       [15:0]   _zz_3073;
  wire       [15:0]   _zz_3074;
  wire       [15:0]   _zz_3075;
  wire       [15:0]   _zz_3076;
  wire       [15:0]   _zz_3077;
  wire       [15:0]   _zz_3078;
  wire       [15:0]   _zz_3079;
  wire       [15:0]   _zz_3080;
  wire       [15:0]   _zz_3081;
  wire       [15:0]   _zz_3082;
  wire       [15:0]   _zz_3083;
  wire       [15:0]   _zz_3084;
  wire       [15:0]   _zz_3085;
  wire       [15:0]   _zz_3086;
  wire       [31:0]   _zz_3087;
  wire       [31:0]   _zz_3088;
  wire       [15:0]   _zz_3089;
  wire       [31:0]   _zz_3090;
  wire       [31:0]   _zz_3091;
  wire       [15:0]   _zz_3092;
  wire       [15:0]   _zz_3093;
  wire       [15:0]   _zz_3094;
  wire       [15:0]   _zz_3095;
  wire       [15:0]   _zz_3096;
  wire       [15:0]   _zz_3097;
  wire       [15:0]   _zz_3098;
  wire       [15:0]   _zz_3099;
  wire       [15:0]   _zz_3100;
  wire       [15:0]   _zz_3101;
  wire       [15:0]   _zz_3102;
  wire       [15:0]   _zz_3103;
  wire       [15:0]   _zz_3104;
  wire       [15:0]   _zz_3105;
  wire       [15:0]   _zz_3106;
  wire       [15:0]   _zz_3107;
  wire       [15:0]   _zz_3108;
  wire       [31:0]   _zz_3109;
  wire       [31:0]   _zz_3110;
  wire       [15:0]   _zz_3111;
  wire       [31:0]   _zz_3112;
  wire       [31:0]   _zz_3113;
  wire       [15:0]   _zz_3114;
  wire       [15:0]   _zz_3115;
  wire       [15:0]   _zz_3116;
  wire       [15:0]   _zz_3117;
  wire       [15:0]   _zz_3118;
  wire       [15:0]   _zz_3119;
  wire       [15:0]   _zz_3120;
  wire       [15:0]   _zz_3121;
  wire       [15:0]   _zz_3122;
  wire       [15:0]   _zz_3123;
  wire       [15:0]   _zz_3124;
  wire       [15:0]   _zz_3125;
  wire       [15:0]   _zz_3126;
  wire       [15:0]   _zz_3127;
  wire       [15:0]   _zz_3128;
  wire       [15:0]   _zz_3129;
  wire       [15:0]   _zz_3130;
  wire       [31:0]   _zz_3131;
  wire       [31:0]   _zz_3132;
  wire       [15:0]   _zz_3133;
  wire       [31:0]   _zz_3134;
  wire       [31:0]   _zz_3135;
  wire       [15:0]   _zz_3136;
  wire       [15:0]   _zz_3137;
  wire       [15:0]   _zz_3138;
  wire       [15:0]   _zz_3139;
  wire       [15:0]   _zz_3140;
  wire       [15:0]   _zz_3141;
  wire       [15:0]   _zz_3142;
  wire       [15:0]   _zz_3143;
  wire       [15:0]   _zz_3144;
  wire       [15:0]   _zz_3145;
  wire       [15:0]   _zz_3146;
  wire       [15:0]   _zz_3147;
  wire       [15:0]   _zz_3148;
  wire       [15:0]   _zz_3149;
  wire       [15:0]   _zz_3150;
  wire       [15:0]   _zz_3151;
  wire       [15:0]   _zz_3152;
  wire       [31:0]   _zz_3153;
  wire       [31:0]   _zz_3154;
  wire       [15:0]   _zz_3155;
  wire       [31:0]   _zz_3156;
  wire       [31:0]   _zz_3157;
  wire       [15:0]   _zz_3158;
  wire       [15:0]   _zz_3159;
  wire       [15:0]   _zz_3160;
  wire       [15:0]   _zz_3161;
  wire       [15:0]   _zz_3162;
  wire       [15:0]   _zz_3163;
  wire       [15:0]   _zz_3164;
  wire       [15:0]   _zz_3165;
  wire       [15:0]   _zz_3166;
  wire       [15:0]   _zz_3167;
  wire       [15:0]   _zz_3168;
  wire       [15:0]   _zz_3169;
  wire       [15:0]   _zz_3170;
  wire       [15:0]   _zz_3171;
  wire       [15:0]   _zz_3172;
  wire       [15:0]   _zz_3173;
  wire       [15:0]   _zz_3174;
  wire       [31:0]   _zz_3175;
  wire       [31:0]   _zz_3176;
  wire       [15:0]   _zz_3177;
  wire       [31:0]   _zz_3178;
  wire       [31:0]   _zz_3179;
  wire       [15:0]   _zz_3180;
  wire       [15:0]   _zz_3181;
  wire       [15:0]   _zz_3182;
  wire       [15:0]   _zz_3183;
  wire       [15:0]   _zz_3184;
  wire       [15:0]   _zz_3185;
  wire       [15:0]   _zz_3186;
  wire       [15:0]   _zz_3187;
  wire       [15:0]   _zz_3188;
  wire       [15:0]   _zz_3189;
  wire       [15:0]   _zz_3190;
  wire       [15:0]   _zz_3191;
  wire       [15:0]   _zz_3192;
  wire       [15:0]   _zz_3193;
  wire       [15:0]   _zz_3194;
  wire       [15:0]   _zz_3195;
  wire       [15:0]   _zz_3196;
  wire       [31:0]   _zz_3197;
  wire       [31:0]   _zz_3198;
  wire       [15:0]   _zz_3199;
  wire       [31:0]   _zz_3200;
  wire       [31:0]   _zz_3201;
  wire       [15:0]   _zz_3202;
  wire       [15:0]   _zz_3203;
  wire       [15:0]   _zz_3204;
  wire       [15:0]   _zz_3205;
  wire       [15:0]   _zz_3206;
  wire       [15:0]   _zz_3207;
  wire       [15:0]   _zz_3208;
  wire       [15:0]   _zz_3209;
  wire       [15:0]   _zz_3210;
  wire       [15:0]   _zz_3211;
  wire       [15:0]   _zz_3212;
  wire       [15:0]   _zz_3213;
  wire       [15:0]   _zz_3214;
  wire       [15:0]   _zz_3215;
  wire       [15:0]   _zz_3216;
  wire       [15:0]   _zz_3217;
  wire       [15:0]   _zz_3218;
  wire       [31:0]   _zz_3219;
  wire       [31:0]   _zz_3220;
  wire       [15:0]   _zz_3221;
  wire       [31:0]   _zz_3222;
  wire       [31:0]   _zz_3223;
  wire       [15:0]   _zz_3224;
  wire       [15:0]   _zz_3225;
  wire       [15:0]   _zz_3226;
  wire       [15:0]   _zz_3227;
  wire       [15:0]   _zz_3228;
  wire       [15:0]   _zz_3229;
  wire       [15:0]   _zz_3230;
  wire       [15:0]   _zz_3231;
  wire       [15:0]   _zz_3232;
  wire       [15:0]   _zz_3233;
  wire       [15:0]   _zz_3234;
  wire       [15:0]   _zz_3235;
  wire       [15:0]   _zz_3236;
  wire       [15:0]   _zz_3237;
  wire       [15:0]   _zz_3238;
  wire       [15:0]   _zz_3239;
  wire       [15:0]   _zz_3240;
  wire       [31:0]   _zz_3241;
  wire       [31:0]   _zz_3242;
  wire       [15:0]   _zz_3243;
  wire       [31:0]   _zz_3244;
  wire       [31:0]   _zz_3245;
  wire       [15:0]   _zz_3246;
  wire       [15:0]   _zz_3247;
  wire       [15:0]   _zz_3248;
  wire       [15:0]   _zz_3249;
  wire       [15:0]   _zz_3250;
  wire       [15:0]   _zz_3251;
  wire       [15:0]   _zz_3252;
  wire       [15:0]   _zz_3253;
  wire       [15:0]   _zz_3254;
  wire       [15:0]   _zz_3255;
  wire       [15:0]   _zz_3256;
  wire       [15:0]   _zz_3257;
  wire       [15:0]   _zz_3258;
  wire       [15:0]   _zz_3259;
  wire       [15:0]   _zz_3260;
  wire       [15:0]   _zz_3261;
  wire       [15:0]   _zz_3262;
  wire       [31:0]   _zz_3263;
  wire       [31:0]   _zz_3264;
  wire       [15:0]   _zz_3265;
  wire       [31:0]   _zz_3266;
  wire       [31:0]   _zz_3267;
  wire       [15:0]   _zz_3268;
  wire       [15:0]   _zz_3269;
  wire       [15:0]   _zz_3270;
  wire       [15:0]   _zz_3271;
  wire       [15:0]   _zz_3272;
  wire       [15:0]   _zz_3273;
  wire       [15:0]   _zz_3274;
  wire       [15:0]   _zz_3275;
  wire       [15:0]   _zz_3276;
  wire       [15:0]   _zz_3277;
  wire       [15:0]   _zz_3278;
  wire       [15:0]   _zz_3279;
  wire       [15:0]   _zz_3280;
  wire       [15:0]   _zz_3281;
  wire       [15:0]   _zz_3282;
  wire       [15:0]   _zz_3283;
  wire       [15:0]   _zz_3284;
  wire       [31:0]   _zz_3285;
  wire       [31:0]   _zz_3286;
  wire       [15:0]   _zz_3287;
  wire       [31:0]   _zz_3288;
  wire       [31:0]   _zz_3289;
  wire       [15:0]   _zz_3290;
  wire       [15:0]   _zz_3291;
  wire       [15:0]   _zz_3292;
  wire       [15:0]   _zz_3293;
  wire       [15:0]   _zz_3294;
  wire       [15:0]   _zz_3295;
  wire       [15:0]   _zz_3296;
  wire       [15:0]   _zz_3297;
  wire       [15:0]   _zz_3298;
  wire       [15:0]   _zz_3299;
  wire       [15:0]   _zz_3300;
  wire       [15:0]   _zz_3301;
  wire       [15:0]   _zz_3302;
  wire       [15:0]   _zz_3303;
  wire       [15:0]   _zz_3304;
  wire       [15:0]   _zz_3305;
  wire       [15:0]   _zz_3306;
  wire       [31:0]   _zz_3307;
  wire       [31:0]   _zz_3308;
  wire       [15:0]   _zz_3309;
  wire       [31:0]   _zz_3310;
  wire       [31:0]   _zz_3311;
  wire       [15:0]   _zz_3312;
  wire       [15:0]   _zz_3313;
  wire       [15:0]   _zz_3314;
  wire       [15:0]   _zz_3315;
  wire       [15:0]   _zz_3316;
  wire       [15:0]   _zz_3317;
  wire       [15:0]   _zz_3318;
  wire       [15:0]   _zz_3319;
  wire       [15:0]   _zz_3320;
  wire       [15:0]   _zz_3321;
  wire       [15:0]   _zz_3322;
  wire       [15:0]   _zz_3323;
  wire       [15:0]   _zz_3324;
  wire       [15:0]   _zz_3325;
  wire       [15:0]   _zz_3326;
  wire       [15:0]   _zz_3327;
  wire       [15:0]   _zz_3328;
  wire       [31:0]   _zz_3329;
  wire       [31:0]   _zz_3330;
  wire       [15:0]   _zz_3331;
  wire       [31:0]   _zz_3332;
  wire       [31:0]   _zz_3333;
  wire       [15:0]   _zz_3334;
  wire       [15:0]   _zz_3335;
  wire       [15:0]   _zz_3336;
  wire       [15:0]   _zz_3337;
  wire       [15:0]   _zz_3338;
  wire       [15:0]   _zz_3339;
  wire       [15:0]   _zz_3340;
  wire       [15:0]   _zz_3341;
  wire       [15:0]   _zz_3342;
  wire       [15:0]   _zz_3343;
  wire       [15:0]   _zz_3344;
  wire       [15:0]   _zz_3345;
  wire       [15:0]   _zz_3346;
  wire       [15:0]   _zz_3347;
  wire       [15:0]   _zz_3348;
  wire       [15:0]   _zz_3349;
  wire       [15:0]   _zz_3350;
  wire       [31:0]   _zz_3351;
  wire       [31:0]   _zz_3352;
  wire       [15:0]   _zz_3353;
  wire       [31:0]   _zz_3354;
  wire       [31:0]   _zz_3355;
  wire       [15:0]   _zz_3356;
  wire       [15:0]   _zz_3357;
  wire       [15:0]   _zz_3358;
  wire       [15:0]   _zz_3359;
  wire       [15:0]   _zz_3360;
  wire       [15:0]   _zz_3361;
  wire       [15:0]   _zz_3362;
  wire       [15:0]   _zz_3363;
  wire       [15:0]   _zz_3364;
  wire       [15:0]   _zz_3365;
  wire       [15:0]   _zz_3366;
  wire       [15:0]   _zz_3367;
  wire       [15:0]   _zz_3368;
  wire       [15:0]   _zz_3369;
  wire       [15:0]   _zz_3370;
  wire       [15:0]   _zz_3371;
  wire       [15:0]   _zz_3372;
  wire       [31:0]   _zz_3373;
  wire       [31:0]   _zz_3374;
  wire       [15:0]   _zz_3375;
  wire       [31:0]   _zz_3376;
  wire       [31:0]   _zz_3377;
  wire       [15:0]   _zz_3378;
  wire       [15:0]   _zz_3379;
  wire       [15:0]   _zz_3380;
  wire       [15:0]   _zz_3381;
  wire       [15:0]   _zz_3382;
  wire       [15:0]   _zz_3383;
  wire       [15:0]   _zz_3384;
  wire       [15:0]   _zz_3385;
  wire       [15:0]   _zz_3386;
  wire       [15:0]   _zz_3387;
  wire       [15:0]   _zz_3388;
  wire       [15:0]   _zz_3389;
  wire       [15:0]   _zz_3390;
  wire       [15:0]   _zz_3391;
  wire       [15:0]   _zz_3392;
  wire       [15:0]   _zz_3393;
  wire       [15:0]   _zz_3394;
  wire       [31:0]   _zz_3395;
  wire       [31:0]   _zz_3396;
  wire       [15:0]   _zz_3397;
  wire       [31:0]   _zz_3398;
  wire       [31:0]   _zz_3399;
  wire       [15:0]   _zz_3400;
  wire       [15:0]   _zz_3401;
  wire       [15:0]   _zz_3402;
  wire       [15:0]   _zz_3403;
  wire       [15:0]   _zz_3404;
  wire       [15:0]   _zz_3405;
  wire       [15:0]   _zz_3406;
  wire       [15:0]   _zz_3407;
  wire       [15:0]   _zz_3408;
  wire       [15:0]   _zz_3409;
  wire       [15:0]   _zz_3410;
  wire       [15:0]   _zz_3411;
  wire       [15:0]   _zz_3412;
  wire       [15:0]   _zz_3413;
  wire       [15:0]   _zz_3414;
  wire       [15:0]   _zz_3415;
  wire       [15:0]   _zz_3416;
  wire       [31:0]   _zz_3417;
  wire       [31:0]   _zz_3418;
  wire       [15:0]   _zz_3419;
  wire       [31:0]   _zz_3420;
  wire       [31:0]   _zz_3421;
  wire       [15:0]   _zz_3422;
  wire       [15:0]   _zz_3423;
  wire       [15:0]   _zz_3424;
  wire       [15:0]   _zz_3425;
  wire       [15:0]   _zz_3426;
  wire       [15:0]   _zz_3427;
  wire       [15:0]   _zz_3428;
  wire       [15:0]   _zz_3429;
  wire       [15:0]   _zz_3430;
  wire       [15:0]   _zz_3431;
  wire       [15:0]   _zz_3432;
  wire       [15:0]   _zz_3433;
  wire       [15:0]   _zz_3434;
  wire       [15:0]   _zz_3435;
  wire       [15:0]   _zz_3436;
  wire       [15:0]   _zz_3437;
  wire       [15:0]   _zz_3438;
  wire       [31:0]   _zz_3439;
  wire       [31:0]   _zz_3440;
  wire       [15:0]   _zz_3441;
  wire       [31:0]   _zz_3442;
  wire       [31:0]   _zz_3443;
  wire       [15:0]   _zz_3444;
  wire       [15:0]   _zz_3445;
  wire       [15:0]   _zz_3446;
  wire       [15:0]   _zz_3447;
  wire       [15:0]   _zz_3448;
  wire       [15:0]   _zz_3449;
  wire       [15:0]   _zz_3450;
  wire       [15:0]   _zz_3451;
  wire       [15:0]   _zz_3452;
  wire       [15:0]   _zz_3453;
  wire       [15:0]   _zz_3454;
  wire       [15:0]   _zz_3455;
  wire       [15:0]   _zz_3456;
  wire       [15:0]   _zz_3457;
  wire       [15:0]   _zz_3458;
  wire       [15:0]   _zz_3459;
  wire       [15:0]   _zz_3460;
  wire       [31:0]   _zz_3461;
  wire       [31:0]   _zz_3462;
  wire       [15:0]   _zz_3463;
  wire       [31:0]   _zz_3464;
  wire       [31:0]   _zz_3465;
  wire       [15:0]   _zz_3466;
  wire       [15:0]   _zz_3467;
  wire       [15:0]   _zz_3468;
  wire       [15:0]   _zz_3469;
  wire       [15:0]   _zz_3470;
  wire       [15:0]   _zz_3471;
  wire       [15:0]   _zz_3472;
  wire       [15:0]   _zz_3473;
  wire       [15:0]   _zz_3474;
  wire       [15:0]   _zz_3475;
  wire       [15:0]   _zz_3476;
  wire       [15:0]   _zz_3477;
  wire       [15:0]   _zz_3478;
  wire       [15:0]   _zz_3479;
  wire       [15:0]   _zz_3480;
  wire       [15:0]   _zz_3481;
  wire       [15:0]   _zz_3482;
  wire       [31:0]   _zz_3483;
  wire       [31:0]   _zz_3484;
  wire       [15:0]   _zz_3485;
  wire       [31:0]   _zz_3486;
  wire       [31:0]   _zz_3487;
  wire       [15:0]   _zz_3488;
  wire       [15:0]   _zz_3489;
  wire       [15:0]   _zz_3490;
  wire       [15:0]   _zz_3491;
  wire       [15:0]   _zz_3492;
  wire       [15:0]   _zz_3493;
  wire       [15:0]   _zz_3494;
  wire       [15:0]   _zz_3495;
  wire       [15:0]   _zz_3496;
  wire       [15:0]   _zz_3497;
  wire       [15:0]   _zz_3498;
  wire       [15:0]   _zz_3499;
  wire       [15:0]   _zz_3500;
  wire       [15:0]   _zz_3501;
  wire       [15:0]   _zz_3502;
  wire       [15:0]   _zz_3503;
  wire       [15:0]   _zz_3504;
  wire       [31:0]   _zz_3505;
  wire       [31:0]   _zz_3506;
  wire       [15:0]   _zz_3507;
  wire       [31:0]   _zz_3508;
  wire       [31:0]   _zz_3509;
  wire       [15:0]   _zz_3510;
  wire       [15:0]   _zz_3511;
  wire       [15:0]   _zz_3512;
  wire       [15:0]   _zz_3513;
  wire       [15:0]   _zz_3514;
  wire       [15:0]   _zz_3515;
  wire       [15:0]   _zz_3516;
  wire       [15:0]   _zz_3517;
  wire       [15:0]   _zz_3518;
  wire       [15:0]   _zz_3519;
  wire       [15:0]   _zz_3520;
  wire       [15:0]   _zz_3521;
  wire       [15:0]   _zz_3522;
  wire       [15:0]   _zz_3523;
  wire       [15:0]   _zz_3524;
  wire       [15:0]   _zz_3525;
  wire       [15:0]   _zz_3526;
  wire       [31:0]   _zz_3527;
  wire       [31:0]   _zz_3528;
  wire       [15:0]   _zz_3529;
  wire       [31:0]   _zz_3530;
  wire       [31:0]   _zz_3531;
  wire       [15:0]   _zz_3532;
  wire       [15:0]   _zz_3533;
  wire       [15:0]   _zz_3534;
  wire       [15:0]   _zz_3535;
  wire       [15:0]   _zz_3536;
  wire       [15:0]   _zz_3537;
  wire       [15:0]   _zz_3538;
  wire       [15:0]   _zz_3539;
  wire       [15:0]   _zz_3540;
  wire       [15:0]   _zz_3541;
  wire       [15:0]   _zz_3542;
  wire       [15:0]   _zz_3543;
  wire       [15:0]   _zz_3544;
  wire       [15:0]   _zz_3545;
  wire       [15:0]   _zz_3546;
  wire       [15:0]   _zz_3547;
  wire       [15:0]   _zz_3548;
  wire       [31:0]   _zz_3549;
  wire       [31:0]   _zz_3550;
  wire       [15:0]   _zz_3551;
  wire       [31:0]   _zz_3552;
  wire       [31:0]   _zz_3553;
  wire       [15:0]   _zz_3554;
  wire       [15:0]   _zz_3555;
  wire       [15:0]   _zz_3556;
  wire       [15:0]   _zz_3557;
  wire       [15:0]   _zz_3558;
  wire       [15:0]   _zz_3559;
  wire       [15:0]   _zz_3560;
  wire       [15:0]   _zz_3561;
  wire       [15:0]   _zz_3562;
  wire       [15:0]   _zz_3563;
  wire       [15:0]   _zz_3564;
  wire       [15:0]   _zz_3565;
  wire       [15:0]   _zz_3566;
  wire       [15:0]   _zz_3567;
  wire       [15:0]   _zz_3568;
  wire       [15:0]   _zz_3569;
  wire       [15:0]   _zz_3570;
  wire       [31:0]   _zz_3571;
  wire       [31:0]   _zz_3572;
  wire       [15:0]   _zz_3573;
  wire       [31:0]   _zz_3574;
  wire       [31:0]   _zz_3575;
  wire       [15:0]   _zz_3576;
  wire       [15:0]   _zz_3577;
  wire       [15:0]   _zz_3578;
  wire       [15:0]   _zz_3579;
  wire       [15:0]   _zz_3580;
  wire       [15:0]   _zz_3581;
  wire       [15:0]   _zz_3582;
  wire       [15:0]   _zz_3583;
  wire       [15:0]   _zz_3584;
  wire       [15:0]   _zz_3585;
  wire       [15:0]   _zz_3586;
  wire       [15:0]   _zz_3587;
  wire       [15:0]   _zz_3588;
  wire       [15:0]   _zz_3589;
  wire       [15:0]   _zz_3590;
  wire       [15:0]   _zz_3591;
  wire       [15:0]   _zz_3592;
  wire       [31:0]   _zz_3593;
  wire       [31:0]   _zz_3594;
  wire       [15:0]   _zz_3595;
  wire       [31:0]   _zz_3596;
  wire       [31:0]   _zz_3597;
  wire       [15:0]   _zz_3598;
  wire       [15:0]   _zz_3599;
  wire       [15:0]   _zz_3600;
  wire       [15:0]   _zz_3601;
  wire       [15:0]   _zz_3602;
  wire       [15:0]   _zz_3603;
  wire       [15:0]   _zz_3604;
  wire       [15:0]   _zz_3605;
  wire       [15:0]   _zz_3606;
  wire       [15:0]   _zz_3607;
  wire       [15:0]   _zz_3608;
  wire       [15:0]   _zz_3609;
  wire       [15:0]   _zz_3610;
  wire       [15:0]   _zz_3611;
  wire       [15:0]   _zz_3612;
  wire       [15:0]   _zz_3613;
  wire       [15:0]   _zz_3614;
  wire       [31:0]   _zz_3615;
  wire       [31:0]   _zz_3616;
  wire       [15:0]   _zz_3617;
  wire       [31:0]   _zz_3618;
  wire       [31:0]   _zz_3619;
  wire       [15:0]   _zz_3620;
  wire       [15:0]   _zz_3621;
  wire       [15:0]   _zz_3622;
  wire       [15:0]   _zz_3623;
  wire       [15:0]   _zz_3624;
  wire       [15:0]   _zz_3625;
  wire       [15:0]   _zz_3626;
  wire       [15:0]   _zz_3627;
  wire       [15:0]   _zz_3628;
  wire       [15:0]   _zz_3629;
  wire       [15:0]   _zz_3630;
  wire       [15:0]   _zz_3631;
  wire       [15:0]   _zz_3632;
  wire       [15:0]   _zz_3633;
  wire       [15:0]   _zz_3634;
  wire       [15:0]   _zz_3635;
  wire       [15:0]   _zz_3636;
  wire       [31:0]   _zz_3637;
  wire       [31:0]   _zz_3638;
  wire       [15:0]   _zz_3639;
  wire       [31:0]   _zz_3640;
  wire       [31:0]   _zz_3641;
  wire       [15:0]   _zz_3642;
  wire       [15:0]   _zz_3643;
  wire       [15:0]   _zz_3644;
  wire       [15:0]   _zz_3645;
  wire       [15:0]   _zz_3646;
  wire       [15:0]   _zz_3647;
  wire       [15:0]   _zz_3648;
  wire       [15:0]   _zz_3649;
  wire       [15:0]   _zz_3650;
  wire       [15:0]   _zz_3651;
  wire       [15:0]   _zz_3652;
  wire       [15:0]   _zz_3653;
  wire       [15:0]   _zz_3654;
  wire       [15:0]   _zz_3655;
  wire       [15:0]   _zz_3656;
  wire       [15:0]   _zz_3657;
  wire       [15:0]   _zz_3658;
  wire       [31:0]   _zz_3659;
  wire       [31:0]   _zz_3660;
  wire       [15:0]   _zz_3661;
  wire       [31:0]   _zz_3662;
  wire       [31:0]   _zz_3663;
  wire       [15:0]   _zz_3664;
  wire       [15:0]   _zz_3665;
  wire       [15:0]   _zz_3666;
  wire       [15:0]   _zz_3667;
  wire       [15:0]   _zz_3668;
  wire       [15:0]   _zz_3669;
  wire       [15:0]   _zz_3670;
  wire       [15:0]   _zz_3671;
  wire       [15:0]   _zz_3672;
  wire       [15:0]   _zz_3673;
  wire       [15:0]   _zz_3674;
  wire       [15:0]   _zz_3675;
  wire       [15:0]   _zz_3676;
  wire       [15:0]   _zz_3677;
  wire       [15:0]   _zz_3678;
  wire       [15:0]   _zz_3679;
  wire       [15:0]   _zz_3680;
  wire       [31:0]   _zz_3681;
  wire       [31:0]   _zz_3682;
  wire       [15:0]   _zz_3683;
  wire       [31:0]   _zz_3684;
  wire       [31:0]   _zz_3685;
  wire       [15:0]   _zz_3686;
  wire       [15:0]   _zz_3687;
  wire       [15:0]   _zz_3688;
  wire       [15:0]   _zz_3689;
  wire       [15:0]   _zz_3690;
  wire       [15:0]   _zz_3691;
  wire       [15:0]   _zz_3692;
  wire       [15:0]   _zz_3693;
  wire       [15:0]   _zz_3694;
  wire       [15:0]   _zz_3695;
  wire       [15:0]   _zz_3696;
  wire       [15:0]   _zz_3697;
  wire       [15:0]   _zz_3698;
  wire       [15:0]   _zz_3699;
  wire       [15:0]   _zz_3700;
  wire       [15:0]   _zz_3701;
  wire       [15:0]   _zz_3702;
  wire       [31:0]   _zz_3703;
  wire       [31:0]   _zz_3704;
  wire       [15:0]   _zz_3705;
  wire       [31:0]   _zz_3706;
  wire       [31:0]   _zz_3707;
  wire       [15:0]   _zz_3708;
  wire       [15:0]   _zz_3709;
  wire       [15:0]   _zz_3710;
  wire       [15:0]   _zz_3711;
  wire       [15:0]   _zz_3712;
  wire       [15:0]   _zz_3713;
  wire       [15:0]   _zz_3714;
  wire       [15:0]   _zz_3715;
  wire       [15:0]   _zz_3716;
  wire       [15:0]   _zz_3717;
  wire       [15:0]   _zz_3718;
  wire       [15:0]   _zz_3719;
  wire       [15:0]   _zz_3720;
  wire       [15:0]   _zz_3721;
  wire       [15:0]   _zz_3722;
  wire       [15:0]   _zz_3723;
  wire       [15:0]   _zz_3724;
  wire       [31:0]   _zz_3725;
  wire       [31:0]   _zz_3726;
  wire       [15:0]   _zz_3727;
  wire       [31:0]   _zz_3728;
  wire       [31:0]   _zz_3729;
  wire       [15:0]   _zz_3730;
  wire       [15:0]   _zz_3731;
  wire       [15:0]   _zz_3732;
  wire       [15:0]   _zz_3733;
  wire       [15:0]   _zz_3734;
  wire       [15:0]   _zz_3735;
  wire       [15:0]   _zz_3736;
  wire       [15:0]   _zz_3737;
  wire       [15:0]   _zz_3738;
  wire       [15:0]   _zz_3739;
  wire       [15:0]   _zz_3740;
  wire       [15:0]   _zz_3741;
  wire       [15:0]   _zz_3742;
  wire       [15:0]   _zz_3743;
  wire       [15:0]   _zz_3744;
  wire       [15:0]   _zz_3745;
  wire       [15:0]   _zz_3746;
  wire       [31:0]   _zz_3747;
  wire       [31:0]   _zz_3748;
  wire       [15:0]   _zz_3749;
  wire       [31:0]   _zz_3750;
  wire       [31:0]   _zz_3751;
  wire       [15:0]   _zz_3752;
  wire       [15:0]   _zz_3753;
  wire       [15:0]   _zz_3754;
  wire       [15:0]   _zz_3755;
  wire       [15:0]   _zz_3756;
  wire       [15:0]   _zz_3757;
  wire       [15:0]   _zz_3758;
  wire       [15:0]   _zz_3759;
  wire       [15:0]   _zz_3760;
  wire       [15:0]   _zz_3761;
  wire       [15:0]   _zz_3762;
  wire       [15:0]   _zz_3763;
  wire       [15:0]   _zz_3764;
  wire       [15:0]   _zz_3765;
  wire       [15:0]   _zz_3766;
  wire       [15:0]   _zz_3767;
  wire       [15:0]   _zz_3768;
  wire       [31:0]   _zz_3769;
  wire       [31:0]   _zz_3770;
  wire       [15:0]   _zz_3771;
  wire       [31:0]   _zz_3772;
  wire       [31:0]   _zz_3773;
  wire       [15:0]   _zz_3774;
  wire       [15:0]   _zz_3775;
  wire       [15:0]   _zz_3776;
  wire       [15:0]   _zz_3777;
  wire       [15:0]   _zz_3778;
  wire       [15:0]   _zz_3779;
  wire       [15:0]   _zz_3780;
  wire       [15:0]   _zz_3781;
  wire       [15:0]   _zz_3782;
  wire       [15:0]   _zz_3783;
  wire       [15:0]   _zz_3784;
  wire       [15:0]   _zz_3785;
  wire       [15:0]   _zz_3786;
  wire       [15:0]   _zz_3787;
  wire       [15:0]   _zz_3788;
  wire       [15:0]   _zz_3789;
  wire       [15:0]   _zz_3790;
  wire       [31:0]   _zz_3791;
  wire       [31:0]   _zz_3792;
  wire       [15:0]   _zz_3793;
  wire       [31:0]   _zz_3794;
  wire       [31:0]   _zz_3795;
  wire       [15:0]   _zz_3796;
  wire       [15:0]   _zz_3797;
  wire       [15:0]   _zz_3798;
  wire       [15:0]   _zz_3799;
  wire       [15:0]   _zz_3800;
  wire       [15:0]   _zz_3801;
  wire       [15:0]   _zz_3802;
  wire       [15:0]   _zz_3803;
  wire       [15:0]   _zz_3804;
  wire       [15:0]   _zz_3805;
  wire       [15:0]   _zz_3806;
  wire       [15:0]   _zz_3807;
  wire       [15:0]   _zz_3808;
  wire       [15:0]   _zz_3809;
  wire       [15:0]   _zz_3810;
  wire       [15:0]   _zz_3811;
  wire       [15:0]   _zz_3812;
  wire       [31:0]   _zz_3813;
  wire       [31:0]   _zz_3814;
  wire       [15:0]   _zz_3815;
  wire       [31:0]   _zz_3816;
  wire       [31:0]   _zz_3817;
  wire       [15:0]   _zz_3818;
  wire       [15:0]   _zz_3819;
  wire       [15:0]   _zz_3820;
  wire       [15:0]   _zz_3821;
  wire       [15:0]   _zz_3822;
  wire       [15:0]   _zz_3823;
  wire       [15:0]   _zz_3824;
  wire       [15:0]   _zz_3825;
  wire       [15:0]   _zz_3826;
  wire       [15:0]   _zz_3827;
  wire       [15:0]   _zz_3828;
  wire       [15:0]   _zz_3829;
  wire       [15:0]   _zz_3830;
  wire       [15:0]   _zz_3831;
  wire       [15:0]   _zz_3832;
  wire       [15:0]   _zz_3833;
  wire       [15:0]   _zz_3834;
  wire       [31:0]   _zz_3835;
  wire       [31:0]   _zz_3836;
  wire       [15:0]   _zz_3837;
  wire       [31:0]   _zz_3838;
  wire       [31:0]   _zz_3839;
  wire       [15:0]   _zz_3840;
  wire       [15:0]   _zz_3841;
  wire       [15:0]   _zz_3842;
  wire       [15:0]   _zz_3843;
  wire       [15:0]   _zz_3844;
  wire       [15:0]   _zz_3845;
  wire       [15:0]   _zz_3846;
  wire       [15:0]   _zz_3847;
  wire       [15:0]   _zz_3848;
  wire       [15:0]   _zz_3849;
  wire       [15:0]   _zz_3850;
  wire       [15:0]   _zz_3851;
  wire       [15:0]   _zz_3852;
  wire       [15:0]   _zz_3853;
  wire       [15:0]   _zz_3854;
  wire       [15:0]   _zz_3855;
  wire       [15:0]   _zz_3856;
  wire       [31:0]   _zz_3857;
  wire       [31:0]   _zz_3858;
  wire       [15:0]   _zz_3859;
  wire       [31:0]   _zz_3860;
  wire       [31:0]   _zz_3861;
  wire       [15:0]   _zz_3862;
  wire       [15:0]   _zz_3863;
  wire       [15:0]   _zz_3864;
  wire       [15:0]   _zz_3865;
  wire       [15:0]   _zz_3866;
  wire       [15:0]   _zz_3867;
  wire       [15:0]   _zz_3868;
  wire       [15:0]   _zz_3869;
  wire       [15:0]   _zz_3870;
  wire       [15:0]   _zz_3871;
  wire       [15:0]   _zz_3872;
  wire       [15:0]   _zz_3873;
  wire       [15:0]   _zz_3874;
  wire       [15:0]   _zz_3875;
  wire       [15:0]   _zz_3876;
  wire       [15:0]   _zz_3877;
  wire       [15:0]   _zz_3878;
  wire       [31:0]   _zz_3879;
  wire       [31:0]   _zz_3880;
  wire       [15:0]   _zz_3881;
  wire       [31:0]   _zz_3882;
  wire       [31:0]   _zz_3883;
  wire       [15:0]   _zz_3884;
  wire       [15:0]   _zz_3885;
  wire       [15:0]   _zz_3886;
  wire       [15:0]   _zz_3887;
  wire       [15:0]   _zz_3888;
  wire       [15:0]   _zz_3889;
  wire       [15:0]   _zz_3890;
  wire       [15:0]   _zz_3891;
  wire       [15:0]   _zz_3892;
  wire       [15:0]   _zz_3893;
  wire       [15:0]   _zz_3894;
  wire       [15:0]   _zz_3895;
  wire       [15:0]   _zz_3896;
  wire       [15:0]   _zz_3897;
  wire       [15:0]   _zz_3898;
  wire       [15:0]   _zz_3899;
  wire       [15:0]   _zz_3900;
  wire       [31:0]   _zz_3901;
  wire       [31:0]   _zz_3902;
  wire       [15:0]   _zz_3903;
  wire       [31:0]   _zz_3904;
  wire       [31:0]   _zz_3905;
  wire       [15:0]   _zz_3906;
  wire       [15:0]   _zz_3907;
  wire       [15:0]   _zz_3908;
  wire       [15:0]   _zz_3909;
  wire       [15:0]   _zz_3910;
  wire       [15:0]   _zz_3911;
  wire       [15:0]   _zz_3912;
  wire       [15:0]   _zz_3913;
  wire       [15:0]   _zz_3914;
  wire       [15:0]   _zz_3915;
  wire       [15:0]   _zz_3916;
  wire       [15:0]   _zz_3917;
  wire       [15:0]   _zz_3918;
  wire       [15:0]   _zz_3919;
  wire       [15:0]   _zz_3920;
  wire       [15:0]   _zz_3921;
  wire       [15:0]   _zz_3922;
  wire       [31:0]   _zz_3923;
  wire       [31:0]   _zz_3924;
  wire       [15:0]   _zz_3925;
  wire       [31:0]   _zz_3926;
  wire       [31:0]   _zz_3927;
  wire       [15:0]   _zz_3928;
  wire       [15:0]   _zz_3929;
  wire       [15:0]   _zz_3930;
  wire       [15:0]   _zz_3931;
  wire       [15:0]   _zz_3932;
  wire       [15:0]   _zz_3933;
  wire       [15:0]   _zz_3934;
  wire       [15:0]   _zz_3935;
  wire       [15:0]   _zz_3936;
  wire       [15:0]   _zz_3937;
  wire       [15:0]   _zz_3938;
  wire       [15:0]   _zz_3939;
  wire       [15:0]   _zz_3940;
  wire       [15:0]   _zz_3941;
  wire       [15:0]   _zz_3942;
  wire       [15:0]   _zz_3943;
  wire       [15:0]   _zz_3944;
  wire       [31:0]   _zz_3945;
  wire       [31:0]   _zz_3946;
  wire       [15:0]   _zz_3947;
  wire       [31:0]   _zz_3948;
  wire       [31:0]   _zz_3949;
  wire       [15:0]   _zz_3950;
  wire       [15:0]   _zz_3951;
  wire       [15:0]   _zz_3952;
  wire       [15:0]   _zz_3953;
  wire       [15:0]   _zz_3954;
  wire       [15:0]   _zz_3955;
  wire       [15:0]   _zz_3956;
  wire       [15:0]   _zz_3957;
  wire       [15:0]   _zz_3958;
  wire       [15:0]   _zz_3959;
  wire       [15:0]   _zz_3960;
  wire       [15:0]   _zz_3961;
  wire       [15:0]   _zz_3962;
  wire       [15:0]   _zz_3963;
  wire       [15:0]   _zz_3964;
  wire       [15:0]   _zz_3965;
  wire       [15:0]   _zz_3966;
  wire       [31:0]   _zz_3967;
  wire       [31:0]   _zz_3968;
  wire       [15:0]   _zz_3969;
  wire       [31:0]   _zz_3970;
  wire       [31:0]   _zz_3971;
  wire       [15:0]   _zz_3972;
  wire       [15:0]   _zz_3973;
  wire       [15:0]   _zz_3974;
  wire       [15:0]   _zz_3975;
  wire       [15:0]   _zz_3976;
  wire       [15:0]   _zz_3977;
  wire       [15:0]   _zz_3978;
  wire       [15:0]   _zz_3979;
  wire       [15:0]   _zz_3980;
  wire       [15:0]   _zz_3981;
  wire       [15:0]   _zz_3982;
  wire       [15:0]   _zz_3983;
  wire       [15:0]   _zz_3984;
  wire       [15:0]   _zz_3985;
  wire       [15:0]   _zz_3986;
  wire       [15:0]   _zz_3987;
  wire       [15:0]   _zz_3988;
  wire       [31:0]   _zz_3989;
  wire       [31:0]   _zz_3990;
  wire       [15:0]   _zz_3991;
  wire       [31:0]   _zz_3992;
  wire       [31:0]   _zz_3993;
  wire       [15:0]   _zz_3994;
  wire       [15:0]   _zz_3995;
  wire       [15:0]   _zz_3996;
  wire       [15:0]   _zz_3997;
  wire       [15:0]   _zz_3998;
  wire       [15:0]   _zz_3999;
  wire       [15:0]   _zz_4000;
  wire       [15:0]   _zz_4001;
  wire       [15:0]   _zz_4002;
  wire       [15:0]   _zz_4003;
  wire       [15:0]   _zz_4004;
  wire       [15:0]   _zz_4005;
  wire       [15:0]   _zz_4006;
  wire       [15:0]   _zz_4007;
  wire       [15:0]   _zz_4008;
  wire       [15:0]   _zz_4009;
  wire       [15:0]   _zz_4010;
  wire       [31:0]   _zz_4011;
  wire       [31:0]   _zz_4012;
  wire       [15:0]   _zz_4013;
  wire       [31:0]   _zz_4014;
  wire       [31:0]   _zz_4015;
  wire       [15:0]   _zz_4016;
  wire       [15:0]   _zz_4017;
  wire       [15:0]   _zz_4018;
  wire       [15:0]   _zz_4019;
  wire       [15:0]   _zz_4020;
  wire       [15:0]   _zz_4021;
  wire       [15:0]   _zz_4022;
  wire       [15:0]   _zz_4023;
  wire       [15:0]   _zz_4024;
  wire       [15:0]   _zz_4025;
  wire       [15:0]   _zz_4026;
  wire       [15:0]   _zz_4027;
  wire       [15:0]   _zz_4028;
  wire       [15:0]   _zz_4029;
  wire       [15:0]   _zz_4030;
  wire       [15:0]   _zz_4031;
  wire       [15:0]   _zz_4032;
  wire       [31:0]   _zz_4033;
  wire       [31:0]   _zz_4034;
  wire       [15:0]   _zz_4035;
  wire       [31:0]   _zz_4036;
  wire       [31:0]   _zz_4037;
  wire       [15:0]   _zz_4038;
  wire       [15:0]   _zz_4039;
  wire       [15:0]   _zz_4040;
  wire       [15:0]   _zz_4041;
  wire       [15:0]   _zz_4042;
  wire       [15:0]   _zz_4043;
  wire       [15:0]   _zz_4044;
  wire       [15:0]   _zz_4045;
  wire       [15:0]   _zz_4046;
  wire       [15:0]   _zz_4047;
  wire       [15:0]   _zz_4048;
  wire       [15:0]   _zz_4049;
  wire       [15:0]   _zz_4050;
  wire       [15:0]   _zz_4051;
  wire       [15:0]   _zz_4052;
  wire       [15:0]   _zz_4053;
  wire       [15:0]   _zz_4054;
  wire       [31:0]   _zz_4055;
  wire       [31:0]   _zz_4056;
  wire       [15:0]   _zz_4057;
  wire       [31:0]   _zz_4058;
  wire       [31:0]   _zz_4059;
  wire       [15:0]   _zz_4060;
  wire       [15:0]   _zz_4061;
  wire       [15:0]   _zz_4062;
  wire       [15:0]   _zz_4063;
  wire       [15:0]   _zz_4064;
  wire       [15:0]   _zz_4065;
  wire       [15:0]   _zz_4066;
  wire       [15:0]   _zz_4067;
  wire       [15:0]   _zz_4068;
  wire       [15:0]   _zz_4069;
  wire       [15:0]   _zz_4070;
  wire       [15:0]   _zz_4071;
  wire       [15:0]   _zz_4072;
  wire       [15:0]   _zz_4073;
  wire       [15:0]   _zz_4074;
  wire       [15:0]   _zz_4075;
  wire       [15:0]   _zz_4076;
  wire       [31:0]   _zz_4077;
  wire       [31:0]   _zz_4078;
  wire       [15:0]   _zz_4079;
  wire       [31:0]   _zz_4080;
  wire       [31:0]   _zz_4081;
  wire       [15:0]   _zz_4082;
  wire       [15:0]   _zz_4083;
  wire       [15:0]   _zz_4084;
  wire       [15:0]   _zz_4085;
  wire       [15:0]   _zz_4086;
  wire       [15:0]   _zz_4087;
  wire       [15:0]   _zz_4088;
  wire       [15:0]   _zz_4089;
  wire       [15:0]   _zz_4090;
  wire       [15:0]   _zz_4091;
  wire       [15:0]   _zz_4092;
  wire       [15:0]   _zz_4093;
  wire       [15:0]   _zz_4094;
  wire       [15:0]   _zz_4095;
  wire       [15:0]   _zz_4096;
  wire       [15:0]   _zz_4097;
  wire       [15:0]   _zz_4098;
  wire       [31:0]   _zz_4099;
  wire       [31:0]   _zz_4100;
  wire       [15:0]   _zz_4101;
  wire       [31:0]   _zz_4102;
  wire       [31:0]   _zz_4103;
  wire       [15:0]   _zz_4104;
  wire       [15:0]   _zz_4105;
  wire       [15:0]   _zz_4106;
  wire       [15:0]   _zz_4107;
  wire       [15:0]   _zz_4108;
  wire       [15:0]   _zz_4109;
  wire       [15:0]   _zz_4110;
  wire       [15:0]   _zz_4111;
  wire       [15:0]   _zz_4112;
  wire       [15:0]   _zz_4113;
  wire       [15:0]   _zz_4114;
  wire       [15:0]   _zz_4115;
  wire       [15:0]   _zz_4116;
  wire       [15:0]   _zz_4117;
  wire       [15:0]   _zz_4118;
  wire       [15:0]   _zz_4119;
  wire       [15:0]   _zz_4120;
  wire       [31:0]   _zz_4121;
  wire       [31:0]   _zz_4122;
  wire       [15:0]   _zz_4123;
  wire       [31:0]   _zz_4124;
  wire       [31:0]   _zz_4125;
  wire       [15:0]   _zz_4126;
  wire       [15:0]   _zz_4127;
  wire       [15:0]   _zz_4128;
  wire       [15:0]   _zz_4129;
  wire       [15:0]   _zz_4130;
  wire       [15:0]   _zz_4131;
  wire       [15:0]   _zz_4132;
  wire       [15:0]   _zz_4133;
  wire       [15:0]   _zz_4134;
  wire       [15:0]   _zz_4135;
  wire       [15:0]   _zz_4136;
  wire       [15:0]   _zz_4137;
  wire       [15:0]   _zz_4138;
  wire       [15:0]   _zz_4139;
  wire       [15:0]   _zz_4140;
  wire       [15:0]   _zz_4141;
  wire       [15:0]   _zz_4142;
  wire       [31:0]   _zz_4143;
  wire       [31:0]   _zz_4144;
  wire       [15:0]   _zz_4145;
  wire       [31:0]   _zz_4146;
  wire       [31:0]   _zz_4147;
  wire       [15:0]   _zz_4148;
  wire       [15:0]   _zz_4149;
  wire       [15:0]   _zz_4150;
  wire       [15:0]   _zz_4151;
  wire       [15:0]   _zz_4152;
  wire       [15:0]   _zz_4153;
  wire       [15:0]   _zz_4154;
  wire       [15:0]   _zz_4155;
  wire       [15:0]   _zz_4156;
  wire       [15:0]   _zz_4157;
  wire       [15:0]   _zz_4158;
  wire       [15:0]   _zz_4159;
  wire       [15:0]   _zz_4160;
  wire       [15:0]   _zz_4161;
  wire       [15:0]   _zz_4162;
  wire       [15:0]   _zz_4163;
  wire       [15:0]   _zz_4164;
  wire       [31:0]   _zz_4165;
  wire       [31:0]   _zz_4166;
  wire       [15:0]   _zz_4167;
  wire       [31:0]   _zz_4168;
  wire       [31:0]   _zz_4169;
  wire       [15:0]   _zz_4170;
  wire       [15:0]   _zz_4171;
  wire       [15:0]   _zz_4172;
  wire       [15:0]   _zz_4173;
  wire       [15:0]   _zz_4174;
  wire       [15:0]   _zz_4175;
  wire       [15:0]   _zz_4176;
  wire       [15:0]   _zz_4177;
  wire       [15:0]   _zz_4178;
  wire       [15:0]   _zz_4179;
  wire       [15:0]   _zz_4180;
  wire       [15:0]   _zz_4181;
  wire       [15:0]   _zz_4182;
  wire       [15:0]   _zz_4183;
  wire       [15:0]   _zz_4184;
  wire       [15:0]   _zz_4185;
  wire       [15:0]   _zz_4186;
  wire       [31:0]   _zz_4187;
  wire       [31:0]   _zz_4188;
  wire       [15:0]   _zz_4189;
  wire       [31:0]   _zz_4190;
  wire       [31:0]   _zz_4191;
  wire       [15:0]   _zz_4192;
  wire       [15:0]   _zz_4193;
  wire       [15:0]   _zz_4194;
  wire       [15:0]   _zz_4195;
  wire       [15:0]   _zz_4196;
  wire       [15:0]   _zz_4197;
  wire       [15:0]   _zz_4198;
  wire       [15:0]   _zz_4199;
  wire       [15:0]   _zz_4200;
  wire       [15:0]   _zz_4201;
  wire       [15:0]   _zz_4202;
  wire       [15:0]   _zz_4203;
  wire       [15:0]   _zz_4204;
  wire       [15:0]   _zz_4205;
  wire       [15:0]   _zz_4206;
  wire       [15:0]   _zz_4207;
  wire       [15:0]   _zz_4208;
  wire       [31:0]   _zz_4209;
  wire       [31:0]   _zz_4210;
  wire       [15:0]   _zz_4211;
  wire       [31:0]   _zz_4212;
  wire       [31:0]   _zz_4213;
  wire       [15:0]   _zz_4214;
  wire       [15:0]   _zz_4215;
  wire       [15:0]   _zz_4216;
  wire       [15:0]   _zz_4217;
  wire       [15:0]   _zz_4218;
  wire       [15:0]   _zz_4219;
  wire       [15:0]   _zz_4220;
  wire       [15:0]   _zz_4221;
  wire       [15:0]   _zz_4222;
  wire       [15:0]   _zz_4223;
  wire       [15:0]   _zz_4224;
  wire       [15:0]   _zz_4225;
  wire       [15:0]   _zz_4226;
  wire       [15:0]   _zz_4227;
  wire       [15:0]   _zz_4228;
  wire       [15:0]   _zz_4229;
  wire       [15:0]   _zz_4230;
  wire       [31:0]   _zz_4231;
  wire       [31:0]   _zz_4232;
  wire       [15:0]   _zz_4233;
  wire       [31:0]   _zz_4234;
  wire       [31:0]   _zz_4235;
  wire       [15:0]   _zz_4236;
  wire       [15:0]   _zz_4237;
  wire       [15:0]   _zz_4238;
  wire       [15:0]   _zz_4239;
  wire       [15:0]   _zz_4240;
  wire       [15:0]   _zz_4241;
  wire       [15:0]   _zz_4242;
  wire       [15:0]   _zz_4243;
  wire       [15:0]   _zz_4244;
  wire       [15:0]   _zz_4245;
  wire       [15:0]   _zz_4246;
  wire       [15:0]   _zz_4247;
  wire       [15:0]   _zz_4248;
  wire       [15:0]   _zz_4249;
  wire       [15:0]   _zz_4250;
  wire       [15:0]   _zz_4251;
  wire       [15:0]   _zz_4252;
  wire       [31:0]   _zz_4253;
  wire       [31:0]   _zz_4254;
  wire       [15:0]   _zz_4255;
  wire       [31:0]   _zz_4256;
  wire       [31:0]   _zz_4257;
  wire       [15:0]   _zz_4258;
  wire       [15:0]   _zz_4259;
  wire       [15:0]   _zz_4260;
  wire       [15:0]   _zz_4261;
  wire       [15:0]   _zz_4262;
  wire       [15:0]   _zz_4263;
  wire       [15:0]   _zz_4264;
  wire       [15:0]   _zz_4265;
  wire       [15:0]   _zz_4266;
  wire       [15:0]   _zz_4267;
  wire       [15:0]   _zz_4268;
  wire       [15:0]   _zz_4269;
  wire       [15:0]   _zz_4270;
  wire       [15:0]   _zz_4271;
  wire       [15:0]   _zz_4272;
  wire       [15:0]   _zz_4273;
  wire       [15:0]   _zz_4274;
  wire       [31:0]   _zz_4275;
  wire       [31:0]   _zz_4276;
  wire       [15:0]   _zz_4277;
  wire       [31:0]   _zz_4278;
  wire       [31:0]   _zz_4279;
  wire       [15:0]   _zz_4280;
  wire       [15:0]   _zz_4281;
  wire       [15:0]   _zz_4282;
  wire       [15:0]   _zz_4283;
  wire       [15:0]   _zz_4284;
  wire       [15:0]   _zz_4285;
  wire       [15:0]   _zz_4286;
  wire       [15:0]   _zz_4287;
  wire       [15:0]   _zz_4288;
  wire       [15:0]   _zz_4289;
  wire       [15:0]   _zz_4290;
  wire       [15:0]   _zz_4291;
  wire       [15:0]   _zz_4292;
  wire       [15:0]   _zz_4293;
  wire       [15:0]   _zz_4294;
  wire       [15:0]   _zz_4295;
  wire       [15:0]   _zz_4296;
  wire       [31:0]   _zz_4297;
  wire       [31:0]   _zz_4298;
  wire       [15:0]   _zz_4299;
  wire       [31:0]   _zz_4300;
  wire       [31:0]   _zz_4301;
  wire       [15:0]   _zz_4302;
  wire       [15:0]   _zz_4303;
  wire       [15:0]   _zz_4304;
  wire       [15:0]   _zz_4305;
  wire       [15:0]   _zz_4306;
  wire       [15:0]   _zz_4307;
  wire       [15:0]   _zz_4308;
  wire       [15:0]   _zz_4309;
  wire       [15:0]   _zz_4310;
  wire       [15:0]   _zz_4311;
  wire       [15:0]   _zz_4312;
  wire       [15:0]   _zz_4313;
  wire       [15:0]   _zz_4314;
  wire       [15:0]   _zz_4315;
  wire       [15:0]   _zz_4316;
  wire       [15:0]   _zz_4317;
  wire       [15:0]   _zz_4318;
  wire       [31:0]   _zz_4319;
  wire       [31:0]   _zz_4320;
  wire       [15:0]   _zz_4321;
  wire       [31:0]   _zz_4322;
  wire       [31:0]   _zz_4323;
  wire       [15:0]   _zz_4324;
  wire       [15:0]   _zz_4325;
  wire       [15:0]   _zz_4326;
  wire       [15:0]   _zz_4327;
  wire       [15:0]   _zz_4328;
  wire       [15:0]   _zz_4329;
  wire       [15:0]   _zz_4330;
  wire       [15:0]   _zz_4331;
  wire       [15:0]   _zz_4332;
  wire       [15:0]   _zz_4333;
  wire       [15:0]   _zz_4334;
  wire       [15:0]   _zz_4335;
  wire       [15:0]   _zz_4336;
  wire       [15:0]   _zz_4337;
  wire       [15:0]   _zz_4338;
  wire       [15:0]   _zz_4339;
  wire       [15:0]   _zz_4340;
  wire       [31:0]   _zz_4341;
  wire       [31:0]   _zz_4342;
  wire       [15:0]   _zz_4343;
  wire       [31:0]   _zz_4344;
  wire       [31:0]   _zz_4345;
  wire       [15:0]   _zz_4346;
  wire       [15:0]   _zz_4347;
  wire       [15:0]   _zz_4348;
  wire       [15:0]   _zz_4349;
  wire       [15:0]   _zz_4350;
  wire       [15:0]   _zz_4351;
  wire       [15:0]   _zz_4352;
  wire       [15:0]   _zz_4353;
  wire       [15:0]   _zz_4354;
  wire       [15:0]   _zz_4355;
  wire       [15:0]   _zz_4356;
  wire       [15:0]   _zz_4357;
  wire       [15:0]   _zz_4358;
  wire       [15:0]   _zz_4359;
  wire       [15:0]   _zz_4360;
  wire       [15:0]   _zz_4361;
  wire       [15:0]   _zz_4362;
  wire       [31:0]   _zz_4363;
  wire       [31:0]   _zz_4364;
  wire       [15:0]   _zz_4365;
  wire       [31:0]   _zz_4366;
  wire       [31:0]   _zz_4367;
  wire       [15:0]   _zz_4368;
  wire       [15:0]   _zz_4369;
  wire       [15:0]   _zz_4370;
  wire       [15:0]   _zz_4371;
  wire       [15:0]   _zz_4372;
  wire       [15:0]   _zz_4373;
  wire       [15:0]   _zz_4374;
  wire       [15:0]   _zz_4375;
  wire       [15:0]   _zz_4376;
  wire       [15:0]   _zz_4377;
  wire       [15:0]   _zz_4378;
  wire       [15:0]   _zz_4379;
  wire       [15:0]   _zz_4380;
  wire       [15:0]   _zz_4381;
  wire       [15:0]   _zz_4382;
  wire       [15:0]   _zz_4383;
  wire       [15:0]   _zz_4384;
  wire       [31:0]   _zz_4385;
  wire       [31:0]   _zz_4386;
  wire       [15:0]   _zz_4387;
  wire       [31:0]   _zz_4388;
  wire       [31:0]   _zz_4389;
  wire       [15:0]   _zz_4390;
  wire       [15:0]   _zz_4391;
  wire       [15:0]   _zz_4392;
  wire       [15:0]   _zz_4393;
  wire       [15:0]   _zz_4394;
  wire       [15:0]   _zz_4395;
  wire       [15:0]   _zz_4396;
  wire       [15:0]   _zz_4397;
  wire       [15:0]   _zz_4398;
  wire       [15:0]   _zz_4399;
  wire       [15:0]   _zz_4400;
  wire       [15:0]   _zz_4401;
  wire       [15:0]   _zz_4402;
  wire       [15:0]   _zz_4403;
  wire       [15:0]   _zz_4404;
  wire       [15:0]   _zz_4405;
  wire       [15:0]   _zz_4406;
  wire       [31:0]   _zz_4407;
  wire       [31:0]   _zz_4408;
  wire       [15:0]   _zz_4409;
  wire       [31:0]   _zz_4410;
  wire       [31:0]   _zz_4411;
  wire       [15:0]   _zz_4412;
  wire       [15:0]   _zz_4413;
  wire       [15:0]   _zz_4414;
  wire       [15:0]   _zz_4415;
  wire       [15:0]   _zz_4416;
  wire       [15:0]   _zz_4417;
  wire       [15:0]   _zz_4418;
  wire       [15:0]   _zz_4419;
  wire       [15:0]   _zz_4420;
  wire       [15:0]   _zz_4421;
  wire       [15:0]   _zz_4422;
  wire       [15:0]   _zz_4423;
  wire       [15:0]   _zz_4424;
  wire       [15:0]   _zz_4425;
  wire       [15:0]   _zz_4426;
  wire       [15:0]   _zz_4427;
  wire       [15:0]   _zz_4428;
  wire       [31:0]   _zz_4429;
  wire       [31:0]   _zz_4430;
  wire       [15:0]   _zz_4431;
  wire       [31:0]   _zz_4432;
  wire       [31:0]   _zz_4433;
  wire       [15:0]   _zz_4434;
  wire       [15:0]   _zz_4435;
  wire       [15:0]   _zz_4436;
  wire       [15:0]   _zz_4437;
  wire       [15:0]   _zz_4438;
  wire       [15:0]   _zz_4439;
  wire       [15:0]   _zz_4440;
  wire       [15:0]   _zz_4441;
  wire       [15:0]   _zz_4442;
  wire       [15:0]   _zz_4443;
  wire       [15:0]   _zz_4444;
  wire       [15:0]   _zz_4445;
  wire       [15:0]   _zz_4446;
  wire       [15:0]   _zz_4447;
  wire       [15:0]   _zz_4448;
  wire       [15:0]   _zz_4449;
  wire       [15:0]   _zz_4450;
  wire       [31:0]   _zz_4451;
  wire       [31:0]   _zz_4452;
  wire       [15:0]   _zz_4453;
  wire       [31:0]   _zz_4454;
  wire       [31:0]   _zz_4455;
  wire       [15:0]   _zz_4456;
  wire       [15:0]   _zz_4457;
  wire       [15:0]   _zz_4458;
  wire       [15:0]   _zz_4459;
  wire       [15:0]   _zz_4460;
  wire       [15:0]   _zz_4461;
  wire       [15:0]   _zz_4462;
  wire       [15:0]   _zz_4463;
  wire       [15:0]   _zz_4464;
  wire       [15:0]   _zz_4465;
  wire       [15:0]   _zz_4466;
  wire       [15:0]   _zz_4467;
  wire       [15:0]   _zz_4468;
  wire       [15:0]   _zz_4469;
  wire       [15:0]   _zz_4470;
  wire       [15:0]   _zz_4471;
  wire       [15:0]   _zz_4472;
  wire       [31:0]   _zz_4473;
  wire       [31:0]   _zz_4474;
  wire       [15:0]   _zz_4475;
  wire       [31:0]   _zz_4476;
  wire       [31:0]   _zz_4477;
  wire       [15:0]   _zz_4478;
  wire       [15:0]   _zz_4479;
  wire       [15:0]   _zz_4480;
  wire       [15:0]   _zz_4481;
  wire       [15:0]   _zz_4482;
  wire       [15:0]   _zz_4483;
  wire       [15:0]   _zz_4484;
  wire       [15:0]   _zz_4485;
  wire       [15:0]   _zz_4486;
  wire       [15:0]   _zz_4487;
  wire       [15:0]   _zz_4488;
  wire       [15:0]   _zz_4489;
  wire       [15:0]   _zz_4490;
  wire       [15:0]   _zz_4491;
  wire       [15:0]   _zz_4492;
  wire       [15:0]   _zz_4493;
  wire       [15:0]   _zz_4494;
  wire       [31:0]   _zz_4495;
  wire       [31:0]   _zz_4496;
  wire       [15:0]   _zz_4497;
  wire       [31:0]   _zz_4498;
  wire       [31:0]   _zz_4499;
  wire       [15:0]   _zz_4500;
  wire       [15:0]   _zz_4501;
  wire       [15:0]   _zz_4502;
  wire       [15:0]   _zz_4503;
  wire       [15:0]   _zz_4504;
  wire       [15:0]   _zz_4505;
  wire       [15:0]   _zz_4506;
  wire       [15:0]   _zz_4507;
  wire       [15:0]   _zz_4508;
  wire       [15:0]   _zz_4509;
  wire       [15:0]   _zz_4510;
  wire       [15:0]   _zz_4511;
  wire       [15:0]   _zz_4512;
  wire       [15:0]   _zz_4513;
  wire       [15:0]   _zz_4514;
  wire       [15:0]   _zz_4515;
  wire       [15:0]   _zz_4516;
  wire       [31:0]   _zz_4517;
  wire       [31:0]   _zz_4518;
  wire       [15:0]   _zz_4519;
  wire       [31:0]   _zz_4520;
  wire       [31:0]   _zz_4521;
  wire       [15:0]   _zz_4522;
  wire       [15:0]   _zz_4523;
  wire       [15:0]   _zz_4524;
  wire       [15:0]   _zz_4525;
  wire       [15:0]   _zz_4526;
  wire       [15:0]   _zz_4527;
  wire       [15:0]   _zz_4528;
  wire       [15:0]   _zz_4529;
  wire       [15:0]   _zz_4530;
  wire       [15:0]   _zz_4531;
  wire       [15:0]   _zz_4532;
  wire       [15:0]   _zz_4533;
  wire       [15:0]   _zz_4534;
  wire       [15:0]   _zz_4535;
  wire       [15:0]   _zz_4536;
  wire       [15:0]   _zz_4537;
  wire       [15:0]   _zz_4538;
  wire       [31:0]   _zz_4539;
  wire       [31:0]   _zz_4540;
  wire       [15:0]   _zz_4541;
  wire       [31:0]   _zz_4542;
  wire       [31:0]   _zz_4543;
  wire       [15:0]   _zz_4544;
  wire       [15:0]   _zz_4545;
  wire       [15:0]   _zz_4546;
  wire       [15:0]   _zz_4547;
  wire       [15:0]   _zz_4548;
  wire       [15:0]   _zz_4549;
  wire       [15:0]   _zz_4550;
  wire       [15:0]   _zz_4551;
  wire       [15:0]   _zz_4552;
  wire       [15:0]   _zz_4553;
  wire       [15:0]   _zz_4554;
  wire       [15:0]   _zz_4555;
  wire       [15:0]   _zz_4556;
  wire       [15:0]   _zz_4557;
  wire       [15:0]   _zz_4558;
  wire       [15:0]   _zz_4559;
  wire       [15:0]   _zz_4560;
  wire       [31:0]   _zz_4561;
  wire       [31:0]   _zz_4562;
  wire       [15:0]   _zz_4563;
  wire       [31:0]   _zz_4564;
  wire       [31:0]   _zz_4565;
  wire       [15:0]   _zz_4566;
  wire       [15:0]   _zz_4567;
  wire       [15:0]   _zz_4568;
  wire       [15:0]   _zz_4569;
  wire       [15:0]   _zz_4570;
  wire       [15:0]   _zz_4571;
  wire       [15:0]   _zz_4572;
  wire       [15:0]   _zz_4573;
  wire       [15:0]   _zz_4574;
  wire       [15:0]   _zz_4575;
  wire       [15:0]   _zz_4576;
  wire       [15:0]   _zz_4577;
  wire       [15:0]   _zz_4578;
  wire       [15:0]   _zz_4579;
  wire       [15:0]   _zz_4580;
  wire       [15:0]   _zz_4581;
  wire       [15:0]   _zz_4582;
  wire       [31:0]   _zz_4583;
  wire       [31:0]   _zz_4584;
  wire       [15:0]   _zz_4585;
  wire       [31:0]   _zz_4586;
  wire       [31:0]   _zz_4587;
  wire       [15:0]   _zz_4588;
  wire       [15:0]   _zz_4589;
  wire       [15:0]   _zz_4590;
  wire       [15:0]   _zz_4591;
  wire       [15:0]   _zz_4592;
  wire       [15:0]   _zz_4593;
  wire       [15:0]   _zz_4594;
  wire       [15:0]   _zz_4595;
  wire       [15:0]   _zz_4596;
  wire       [15:0]   _zz_4597;
  wire       [15:0]   _zz_4598;
  wire       [15:0]   _zz_4599;
  wire       [15:0]   _zz_4600;
  wire       [15:0]   _zz_4601;
  wire       [15:0]   _zz_4602;
  wire       [15:0]   _zz_4603;
  wire       [15:0]   _zz_4604;
  wire       [31:0]   _zz_4605;
  wire       [31:0]   _zz_4606;
  wire       [15:0]   _zz_4607;
  wire       [31:0]   _zz_4608;
  wire       [31:0]   _zz_4609;
  wire       [15:0]   _zz_4610;
  wire       [15:0]   _zz_4611;
  wire       [15:0]   _zz_4612;
  wire       [15:0]   _zz_4613;
  wire       [15:0]   _zz_4614;
  wire       [15:0]   _zz_4615;
  wire       [15:0]   _zz_4616;
  wire       [15:0]   _zz_4617;
  wire       [15:0]   _zz_4618;
  wire       [15:0]   _zz_4619;
  wire       [15:0]   _zz_4620;
  wire       [15:0]   _zz_4621;
  wire       [15:0]   _zz_4622;
  wire       [15:0]   _zz_4623;
  wire       [15:0]   _zz_4624;
  wire       [15:0]   _zz_4625;
  wire       [15:0]   _zz_4626;
  wire       [31:0]   _zz_4627;
  wire       [31:0]   _zz_4628;
  wire       [15:0]   _zz_4629;
  wire       [31:0]   _zz_4630;
  wire       [31:0]   _zz_4631;
  wire       [15:0]   _zz_4632;
  wire       [15:0]   _zz_4633;
  wire       [15:0]   _zz_4634;
  wire       [15:0]   _zz_4635;
  wire       [15:0]   _zz_4636;
  wire       [15:0]   _zz_4637;
  wire       [15:0]   _zz_4638;
  wire       [15:0]   _zz_4639;
  wire       [15:0]   _zz_4640;
  wire       [15:0]   _zz_4641;
  wire       [15:0]   _zz_4642;
  wire       [15:0]   _zz_4643;
  wire       [15:0]   _zz_4644;
  wire       [15:0]   _zz_4645;
  wire       [15:0]   _zz_4646;
  wire       [15:0]   _zz_4647;
  wire       [15:0]   _zz_4648;
  wire       [31:0]   _zz_4649;
  wire       [31:0]   _zz_4650;
  wire       [15:0]   _zz_4651;
  wire       [31:0]   _zz_4652;
  wire       [31:0]   _zz_4653;
  wire       [15:0]   _zz_4654;
  wire       [15:0]   _zz_4655;
  wire       [15:0]   _zz_4656;
  wire       [15:0]   _zz_4657;
  wire       [15:0]   _zz_4658;
  wire       [15:0]   _zz_4659;
  wire       [15:0]   _zz_4660;
  wire       [15:0]   _zz_4661;
  wire       [15:0]   _zz_4662;
  wire       [15:0]   _zz_4663;
  wire       [15:0]   _zz_4664;
  wire       [15:0]   _zz_4665;
  wire       [15:0]   _zz_4666;
  wire       [15:0]   _zz_4667;
  wire       [15:0]   _zz_4668;
  wire       [15:0]   _zz_4669;
  wire       [15:0]   _zz_4670;
  wire       [31:0]   _zz_4671;
  wire       [31:0]   _zz_4672;
  wire       [15:0]   _zz_4673;
  wire       [31:0]   _zz_4674;
  wire       [31:0]   _zz_4675;
  wire       [15:0]   _zz_4676;
  wire       [15:0]   _zz_4677;
  wire       [15:0]   _zz_4678;
  wire       [15:0]   _zz_4679;
  wire       [15:0]   _zz_4680;
  wire       [15:0]   _zz_4681;
  wire       [15:0]   _zz_4682;
  wire       [15:0]   _zz_4683;
  wire       [15:0]   _zz_4684;
  wire       [15:0]   _zz_4685;
  wire       [15:0]   _zz_4686;
  wire       [15:0]   _zz_4687;
  wire       [15:0]   _zz_4688;
  wire       [15:0]   _zz_4689;
  wire       [15:0]   _zz_4690;
  wire       [15:0]   _zz_4691;
  wire       [15:0]   _zz_4692;
  wire       [31:0]   _zz_4693;
  wire       [31:0]   _zz_4694;
  wire       [15:0]   _zz_4695;
  wire       [31:0]   _zz_4696;
  wire       [31:0]   _zz_4697;
  wire       [15:0]   _zz_4698;
  wire       [15:0]   _zz_4699;
  wire       [15:0]   _zz_4700;
  wire       [15:0]   _zz_4701;
  wire       [15:0]   _zz_4702;
  wire       [15:0]   _zz_4703;
  wire       [15:0]   _zz_4704;
  wire       [15:0]   _zz_4705;
  wire       [15:0]   _zz_4706;
  wire       [15:0]   _zz_4707;
  wire       [15:0]   _zz_4708;
  wire       [15:0]   _zz_4709;
  wire       [15:0]   _zz_4710;
  wire       [15:0]   _zz_4711;
  wire       [15:0]   _zz_4712;
  wire       [15:0]   _zz_4713;
  wire       [15:0]   _zz_4714;
  wire       [31:0]   _zz_4715;
  wire       [31:0]   _zz_4716;
  wire       [15:0]   _zz_4717;
  wire       [31:0]   _zz_4718;
  wire       [31:0]   _zz_4719;
  wire       [15:0]   _zz_4720;
  wire       [15:0]   _zz_4721;
  wire       [15:0]   _zz_4722;
  wire       [15:0]   _zz_4723;
  wire       [15:0]   _zz_4724;
  wire       [15:0]   _zz_4725;
  wire       [15:0]   _zz_4726;
  wire       [15:0]   _zz_4727;
  wire       [15:0]   _zz_4728;
  wire       [15:0]   _zz_4729;
  wire       [15:0]   _zz_4730;
  wire       [15:0]   _zz_4731;
  wire       [15:0]   _zz_4732;
  wire       [15:0]   _zz_4733;
  wire       [15:0]   _zz_4734;
  wire       [15:0]   _zz_4735;
  wire       [15:0]   _zz_4736;
  wire       [31:0]   _zz_4737;
  wire       [31:0]   _zz_4738;
  wire       [15:0]   _zz_4739;
  wire       [31:0]   _zz_4740;
  wire       [31:0]   _zz_4741;
  wire       [15:0]   _zz_4742;
  wire       [15:0]   _zz_4743;
  wire       [15:0]   _zz_4744;
  wire       [15:0]   _zz_4745;
  wire       [15:0]   _zz_4746;
  wire       [15:0]   _zz_4747;
  wire       [15:0]   _zz_4748;
  wire       [15:0]   _zz_4749;
  wire       [15:0]   _zz_4750;
  wire       [15:0]   _zz_4751;
  wire       [15:0]   _zz_4752;
  wire       [15:0]   _zz_4753;
  wire       [15:0]   _zz_4754;
  wire       [15:0]   _zz_4755;
  wire       [15:0]   _zz_4756;
  wire       [15:0]   _zz_4757;
  wire       [15:0]   _zz_4758;
  wire       [31:0]   _zz_4759;
  wire       [31:0]   _zz_4760;
  wire       [15:0]   _zz_4761;
  wire       [31:0]   _zz_4762;
  wire       [31:0]   _zz_4763;
  wire       [15:0]   _zz_4764;
  wire       [15:0]   _zz_4765;
  wire       [15:0]   _zz_4766;
  wire       [15:0]   _zz_4767;
  wire       [15:0]   _zz_4768;
  wire       [15:0]   _zz_4769;
  wire       [15:0]   _zz_4770;
  wire       [15:0]   _zz_4771;
  wire       [15:0]   _zz_4772;
  wire       [15:0]   _zz_4773;
  wire       [15:0]   _zz_4774;
  wire       [15:0]   _zz_4775;
  wire       [15:0]   _zz_4776;
  wire       [15:0]   _zz_4777;
  wire       [15:0]   _zz_4778;
  wire       [15:0]   _zz_4779;
  wire       [15:0]   _zz_4780;
  wire       [31:0]   _zz_4781;
  wire       [31:0]   _zz_4782;
  wire       [15:0]   _zz_4783;
  wire       [31:0]   _zz_4784;
  wire       [31:0]   _zz_4785;
  wire       [15:0]   _zz_4786;
  wire       [15:0]   _zz_4787;
  wire       [15:0]   _zz_4788;
  wire       [15:0]   _zz_4789;
  wire       [15:0]   _zz_4790;
  wire       [15:0]   _zz_4791;
  wire       [15:0]   _zz_4792;
  wire       [15:0]   _zz_4793;
  wire       [15:0]   _zz_4794;
  wire       [15:0]   _zz_4795;
  wire       [15:0]   _zz_4796;
  wire       [15:0]   _zz_4797;
  wire       [15:0]   _zz_4798;
  wire       [15:0]   _zz_4799;
  wire       [15:0]   _zz_4800;
  wire       [15:0]   _zz_4801;
  wire       [15:0]   _zz_4802;
  wire       [31:0]   _zz_4803;
  wire       [31:0]   _zz_4804;
  wire       [15:0]   _zz_4805;
  wire       [31:0]   _zz_4806;
  wire       [31:0]   _zz_4807;
  wire       [15:0]   _zz_4808;
  wire       [15:0]   _zz_4809;
  wire       [15:0]   _zz_4810;
  wire       [15:0]   _zz_4811;
  wire       [15:0]   _zz_4812;
  wire       [15:0]   _zz_4813;
  wire       [15:0]   _zz_4814;
  wire       [15:0]   _zz_4815;
  wire       [15:0]   _zz_4816;
  wire       [15:0]   _zz_4817;
  wire       [15:0]   _zz_4818;
  wire       [15:0]   _zz_4819;
  wire       [15:0]   _zz_4820;
  wire       [15:0]   _zz_4821;
  wire       [15:0]   _zz_4822;
  wire       [15:0]   _zz_4823;
  wire       [15:0]   _zz_4824;
  wire       [31:0]   _zz_4825;
  wire       [31:0]   _zz_4826;
  wire       [15:0]   _zz_4827;
  wire       [31:0]   _zz_4828;
  wire       [31:0]   _zz_4829;
  wire       [15:0]   _zz_4830;
  wire       [15:0]   _zz_4831;
  wire       [15:0]   _zz_4832;
  wire       [15:0]   _zz_4833;
  wire       [15:0]   _zz_4834;
  wire       [15:0]   _zz_4835;
  wire       [15:0]   _zz_4836;
  wire       [15:0]   _zz_4837;
  wire       [15:0]   _zz_4838;
  wire       [15:0]   _zz_4839;
  wire       [15:0]   _zz_4840;
  wire       [15:0]   _zz_4841;
  wire       [15:0]   _zz_4842;
  wire       [15:0]   _zz_4843;
  wire       [15:0]   _zz_4844;
  wire       [15:0]   _zz_4845;
  wire       [15:0]   _zz_4846;
  wire       [31:0]   _zz_4847;
  wire       [31:0]   _zz_4848;
  wire       [15:0]   _zz_4849;
  wire       [31:0]   _zz_4850;
  wire       [31:0]   _zz_4851;
  wire       [15:0]   _zz_4852;
  wire       [15:0]   _zz_4853;
  wire       [15:0]   _zz_4854;
  wire       [15:0]   _zz_4855;
  wire       [15:0]   _zz_4856;
  wire       [15:0]   _zz_4857;
  wire       [15:0]   _zz_4858;
  wire       [15:0]   _zz_4859;
  wire       [15:0]   _zz_4860;
  wire       [15:0]   _zz_4861;
  wire       [15:0]   _zz_4862;
  wire       [15:0]   _zz_4863;
  wire       [15:0]   _zz_4864;
  wire       [15:0]   _zz_4865;
  wire       [15:0]   _zz_4866;
  wire       [15:0]   _zz_4867;
  wire       [15:0]   _zz_4868;
  wire       [31:0]   _zz_4869;
  wire       [31:0]   _zz_4870;
  wire       [15:0]   _zz_4871;
  wire       [31:0]   _zz_4872;
  wire       [31:0]   _zz_4873;
  wire       [15:0]   _zz_4874;
  wire       [15:0]   _zz_4875;
  wire       [15:0]   _zz_4876;
  wire       [15:0]   _zz_4877;
  wire       [15:0]   _zz_4878;
  wire       [15:0]   _zz_4879;
  wire       [15:0]   _zz_4880;
  wire       [15:0]   _zz_4881;
  wire       [15:0]   _zz_4882;
  wire       [15:0]   _zz_4883;
  wire       [15:0]   _zz_4884;
  wire       [15:0]   _zz_4885;
  wire       [15:0]   _zz_4886;
  wire       [15:0]   _zz_4887;
  wire       [15:0]   _zz_4888;
  wire       [15:0]   _zz_4889;
  wire       [15:0]   _zz_4890;
  wire       [31:0]   _zz_4891;
  wire       [31:0]   _zz_4892;
  wire       [15:0]   _zz_4893;
  wire       [31:0]   _zz_4894;
  wire       [31:0]   _zz_4895;
  wire       [15:0]   _zz_4896;
  wire       [15:0]   _zz_4897;
  wire       [15:0]   _zz_4898;
  wire       [15:0]   _zz_4899;
  wire       [15:0]   _zz_4900;
  wire       [15:0]   _zz_4901;
  wire       [15:0]   _zz_4902;
  wire       [15:0]   _zz_4903;
  wire       [15:0]   _zz_4904;
  wire       [15:0]   _zz_4905;
  wire       [15:0]   _zz_4906;
  wire       [15:0]   _zz_4907;
  wire       [15:0]   _zz_4908;
  wire       [15:0]   _zz_4909;
  wire       [15:0]   _zz_4910;
  wire       [15:0]   _zz_4911;
  wire       [15:0]   _zz_4912;
  wire       [31:0]   _zz_4913;
  wire       [31:0]   _zz_4914;
  wire       [15:0]   _zz_4915;
  wire       [31:0]   _zz_4916;
  wire       [31:0]   _zz_4917;
  wire       [15:0]   _zz_4918;
  wire       [15:0]   _zz_4919;
  wire       [15:0]   _zz_4920;
  wire       [15:0]   _zz_4921;
  wire       [15:0]   _zz_4922;
  wire       [15:0]   _zz_4923;
  wire       [15:0]   _zz_4924;
  wire       [15:0]   _zz_4925;
  wire       [15:0]   _zz_4926;
  wire       [15:0]   _zz_4927;
  wire       [15:0]   _zz_4928;
  wire       [15:0]   _zz_4929;
  wire       [15:0]   _zz_4930;
  wire       [15:0]   _zz_4931;
  wire       [15:0]   _zz_4932;
  wire       [15:0]   _zz_4933;
  wire       [15:0]   _zz_4934;
  wire       [31:0]   _zz_4935;
  wire       [31:0]   _zz_4936;
  wire       [15:0]   _zz_4937;
  wire       [31:0]   _zz_4938;
  wire       [31:0]   _zz_4939;
  wire       [15:0]   _zz_4940;
  wire       [15:0]   _zz_4941;
  wire       [15:0]   _zz_4942;
  wire       [15:0]   _zz_4943;
  wire       [15:0]   _zz_4944;
  wire       [15:0]   _zz_4945;
  wire       [15:0]   _zz_4946;
  wire       [15:0]   _zz_4947;
  wire       [15:0]   _zz_4948;
  wire       [15:0]   _zz_4949;
  wire       [15:0]   _zz_4950;
  wire       [15:0]   _zz_4951;
  wire       [15:0]   _zz_4952;
  wire       [15:0]   _zz_4953;
  wire       [15:0]   _zz_4954;
  wire       [15:0]   _zz_4955;
  wire       [15:0]   _zz_4956;
  wire       [31:0]   _zz_4957;
  wire       [31:0]   _zz_4958;
  wire       [15:0]   _zz_4959;
  wire       [31:0]   _zz_4960;
  wire       [31:0]   _zz_4961;
  wire       [15:0]   _zz_4962;
  wire       [15:0]   _zz_4963;
  wire       [15:0]   _zz_4964;
  wire       [15:0]   _zz_4965;
  wire       [15:0]   _zz_4966;
  wire       [15:0]   _zz_4967;
  wire       [15:0]   _zz_4968;
  wire       [15:0]   _zz_4969;
  wire       [15:0]   _zz_4970;
  wire       [15:0]   _zz_4971;
  wire       [15:0]   _zz_4972;
  wire       [15:0]   _zz_4973;
  wire       [15:0]   _zz_4974;
  wire       [15:0]   _zz_4975;
  wire       [15:0]   _zz_4976;
  wire       [15:0]   _zz_4977;
  wire       [15:0]   _zz_4978;
  wire       [31:0]   _zz_4979;
  wire       [31:0]   _zz_4980;
  wire       [15:0]   _zz_4981;
  wire       [31:0]   _zz_4982;
  wire       [31:0]   _zz_4983;
  wire       [15:0]   _zz_4984;
  wire       [15:0]   _zz_4985;
  wire       [15:0]   _zz_4986;
  wire       [15:0]   _zz_4987;
  wire       [15:0]   _zz_4988;
  wire       [15:0]   _zz_4989;
  wire       [15:0]   _zz_4990;
  wire       [15:0]   _zz_4991;
  wire       [15:0]   _zz_4992;
  wire       [15:0]   _zz_4993;
  wire       [15:0]   _zz_4994;
  wire       [15:0]   _zz_4995;
  wire       [15:0]   _zz_4996;
  wire       [15:0]   _zz_4997;
  wire       [15:0]   _zz_4998;
  wire       [15:0]   _zz_4999;
  wire       [15:0]   _zz_5000;
  wire       [31:0]   _zz_5001;
  wire       [31:0]   _zz_5002;
  wire       [15:0]   _zz_5003;
  wire       [31:0]   _zz_5004;
  wire       [31:0]   _zz_5005;
  wire       [15:0]   _zz_5006;
  wire       [15:0]   _zz_5007;
  wire       [15:0]   _zz_5008;
  wire       [15:0]   _zz_5009;
  wire       [15:0]   _zz_5010;
  wire       [15:0]   _zz_5011;
  wire       [15:0]   _zz_5012;
  wire       [15:0]   _zz_5013;
  wire       [15:0]   _zz_5014;
  wire       [15:0]   _zz_5015;
  wire       [15:0]   _zz_5016;
  wire       [15:0]   _zz_5017;
  wire       [15:0]   _zz_5018;
  wire       [15:0]   _zz_5019;
  wire       [15:0]   _zz_5020;
  wire       [15:0]   _zz_5021;
  wire       [15:0]   _zz_5022;
  wire       [31:0]   _zz_5023;
  wire       [31:0]   _zz_5024;
  wire       [15:0]   _zz_5025;
  wire       [31:0]   _zz_5026;
  wire       [31:0]   _zz_5027;
  wire       [15:0]   _zz_5028;
  wire       [15:0]   _zz_5029;
  wire       [15:0]   _zz_5030;
  wire       [15:0]   _zz_5031;
  wire       [15:0]   _zz_5032;
  wire       [15:0]   _zz_5033;
  wire       [15:0]   _zz_5034;
  wire       [15:0]   _zz_5035;
  wire       [15:0]   _zz_5036;
  wire       [15:0]   _zz_5037;
  wire       [15:0]   _zz_5038;
  wire       [15:0]   _zz_5039;
  wire       [15:0]   _zz_5040;
  wire       [15:0]   _zz_5041;
  wire       [15:0]   _zz_5042;
  wire       [15:0]   _zz_5043;
  wire       [15:0]   _zz_5044;
  wire       [31:0]   _zz_5045;
  wire       [31:0]   _zz_5046;
  wire       [15:0]   _zz_5047;
  wire       [31:0]   _zz_5048;
  wire       [31:0]   _zz_5049;
  wire       [15:0]   _zz_5050;
  wire       [15:0]   _zz_5051;
  wire       [15:0]   _zz_5052;
  wire       [15:0]   _zz_5053;
  wire       [15:0]   _zz_5054;
  wire       [15:0]   _zz_5055;
  wire       [15:0]   _zz_5056;
  wire       [15:0]   _zz_5057;
  wire       [15:0]   _zz_5058;
  wire       [15:0]   _zz_5059;
  wire       [15:0]   _zz_5060;
  wire       [15:0]   _zz_5061;
  wire       [15:0]   _zz_5062;
  wire       [15:0]   _zz_5063;
  wire       [15:0]   _zz_5064;
  wire       [15:0]   _zz_5065;
  wire       [15:0]   _zz_5066;
  wire       [31:0]   _zz_5067;
  wire       [31:0]   _zz_5068;
  wire       [15:0]   _zz_5069;
  wire       [31:0]   _zz_5070;
  wire       [31:0]   _zz_5071;
  wire       [15:0]   _zz_5072;
  wire       [15:0]   _zz_5073;
  wire       [15:0]   _zz_5074;
  wire       [15:0]   _zz_5075;
  wire       [15:0]   _zz_5076;
  wire       [15:0]   _zz_5077;
  wire       [15:0]   _zz_5078;
  wire       [15:0]   _zz_5079;
  wire       [15:0]   _zz_5080;
  wire       [15:0]   _zz_5081;
  wire       [15:0]   _zz_5082;
  wire       [15:0]   _zz_5083;
  wire       [15:0]   _zz_5084;
  wire       [15:0]   _zz_5085;
  wire       [15:0]   _zz_5086;
  wire       [15:0]   _zz_5087;
  wire       [15:0]   _zz_5088;
  wire       [31:0]   _zz_5089;
  wire       [31:0]   _zz_5090;
  wire       [15:0]   _zz_5091;
  wire       [31:0]   _zz_5092;
  wire       [31:0]   _zz_5093;
  wire       [15:0]   _zz_5094;
  wire       [15:0]   _zz_5095;
  wire       [15:0]   _zz_5096;
  wire       [15:0]   _zz_5097;
  wire       [15:0]   _zz_5098;
  wire       [15:0]   _zz_5099;
  wire       [15:0]   _zz_5100;
  wire       [15:0]   _zz_5101;
  wire       [15:0]   _zz_5102;
  wire       [15:0]   _zz_5103;
  wire       [15:0]   _zz_5104;
  wire       [15:0]   _zz_5105;
  wire       [15:0]   _zz_5106;
  wire       [15:0]   _zz_5107;
  wire       [15:0]   _zz_5108;
  wire       [15:0]   _zz_5109;
  wire       [15:0]   _zz_5110;
  wire       [31:0]   _zz_5111;
  wire       [31:0]   _zz_5112;
  wire       [15:0]   _zz_5113;
  wire       [31:0]   _zz_5114;
  wire       [31:0]   _zz_5115;
  wire       [15:0]   _zz_5116;
  wire       [15:0]   _zz_5117;
  wire       [15:0]   _zz_5118;
  wire       [15:0]   _zz_5119;
  wire       [15:0]   _zz_5120;
  wire       [15:0]   _zz_5121;
  wire       [15:0]   _zz_5122;
  wire       [15:0]   _zz_5123;
  wire       [15:0]   _zz_5124;
  wire       [15:0]   _zz_5125;
  wire       [15:0]   _zz_5126;
  wire       [15:0]   _zz_5127;
  wire       [15:0]   _zz_5128;
  wire       [15:0]   _zz_5129;
  wire       [15:0]   _zz_5130;
  wire       [15:0]   _zz_5131;
  wire       [15:0]   _zz_5132;
  wire       [31:0]   _zz_5133;
  wire       [31:0]   _zz_5134;
  wire       [15:0]   _zz_5135;
  wire       [31:0]   _zz_5136;
  wire       [31:0]   _zz_5137;
  wire       [15:0]   _zz_5138;
  wire       [15:0]   _zz_5139;
  wire       [15:0]   _zz_5140;
  wire       [15:0]   _zz_5141;
  wire       [15:0]   _zz_5142;
  wire       [15:0]   _zz_5143;
  wire       [15:0]   _zz_5144;
  wire       [15:0]   _zz_5145;
  wire       [15:0]   _zz_5146;
  wire       [15:0]   _zz_5147;
  wire       [15:0]   _zz_5148;
  wire       [15:0]   _zz_5149;
  wire       [15:0]   _zz_5150;
  wire       [15:0]   _zz_5151;
  wire       [15:0]   _zz_5152;
  wire       [15:0]   _zz_5153;
  wire       [15:0]   _zz_5154;
  wire       [31:0]   _zz_5155;
  wire       [31:0]   _zz_5156;
  wire       [15:0]   _zz_5157;
  wire       [31:0]   _zz_5158;
  wire       [31:0]   _zz_5159;
  wire       [15:0]   _zz_5160;
  wire       [15:0]   _zz_5161;
  wire       [15:0]   _zz_5162;
  wire       [15:0]   _zz_5163;
  wire       [15:0]   _zz_5164;
  wire       [15:0]   _zz_5165;
  wire       [15:0]   _zz_5166;
  wire       [15:0]   _zz_5167;
  wire       [15:0]   _zz_5168;
  wire       [15:0]   _zz_5169;
  wire       [15:0]   _zz_5170;
  wire       [15:0]   _zz_5171;
  wire       [15:0]   _zz_5172;
  wire       [15:0]   _zz_5173;
  wire       [15:0]   _zz_5174;
  wire       [15:0]   _zz_5175;
  wire       [15:0]   _zz_5176;
  wire       [31:0]   _zz_5177;
  wire       [31:0]   _zz_5178;
  wire       [15:0]   _zz_5179;
  wire       [31:0]   _zz_5180;
  wire       [31:0]   _zz_5181;
  wire       [15:0]   _zz_5182;
  wire       [15:0]   _zz_5183;
  wire       [15:0]   _zz_5184;
  wire       [15:0]   _zz_5185;
  wire       [15:0]   _zz_5186;
  wire       [15:0]   _zz_5187;
  wire       [15:0]   _zz_5188;
  wire       [15:0]   _zz_5189;
  wire       [15:0]   _zz_5190;
  wire       [15:0]   _zz_5191;
  wire       [15:0]   _zz_5192;
  wire       [15:0]   _zz_5193;
  wire       [15:0]   _zz_5194;
  wire       [15:0]   _zz_5195;
  wire       [15:0]   _zz_5196;
  wire       [15:0]   _zz_5197;
  wire       [15:0]   _zz_5198;
  wire       [31:0]   _zz_5199;
  wire       [31:0]   _zz_5200;
  wire       [15:0]   _zz_5201;
  wire       [31:0]   _zz_5202;
  wire       [31:0]   _zz_5203;
  wire       [15:0]   _zz_5204;
  wire       [15:0]   _zz_5205;
  wire       [15:0]   _zz_5206;
  wire       [15:0]   _zz_5207;
  wire       [15:0]   _zz_5208;
  wire       [15:0]   _zz_5209;
  wire       [15:0]   _zz_5210;
  wire       [15:0]   _zz_5211;
  wire       [15:0]   _zz_5212;
  wire       [15:0]   _zz_5213;
  wire       [15:0]   _zz_5214;
  wire       [15:0]   _zz_5215;
  wire       [15:0]   _zz_5216;
  wire       [15:0]   _zz_5217;
  wire       [15:0]   _zz_5218;
  wire       [15:0]   _zz_5219;
  wire       [15:0]   _zz_5220;
  wire       [31:0]   _zz_5221;
  wire       [31:0]   _zz_5222;
  wire       [15:0]   _zz_5223;
  wire       [31:0]   _zz_5224;
  wire       [31:0]   _zz_5225;
  wire       [15:0]   _zz_5226;
  wire       [15:0]   _zz_5227;
  wire       [15:0]   _zz_5228;
  wire       [15:0]   _zz_5229;
  wire       [15:0]   _zz_5230;
  wire       [15:0]   _zz_5231;
  wire       [15:0]   _zz_5232;
  wire       [15:0]   _zz_5233;
  wire       [15:0]   _zz_5234;
  wire       [15:0]   _zz_5235;
  wire       [15:0]   _zz_5236;
  wire       [15:0]   _zz_5237;
  wire       [15:0]   _zz_5238;
  wire       [15:0]   _zz_5239;
  wire       [15:0]   _zz_5240;
  wire       [15:0]   _zz_5241;
  wire       [15:0]   _zz_5242;
  wire       [31:0]   _zz_5243;
  wire       [31:0]   _zz_5244;
  wire       [15:0]   _zz_5245;
  wire       [31:0]   _zz_5246;
  wire       [31:0]   _zz_5247;
  wire       [15:0]   _zz_5248;
  wire       [15:0]   _zz_5249;
  wire       [15:0]   _zz_5250;
  wire       [15:0]   _zz_5251;
  wire       [15:0]   _zz_5252;
  wire       [15:0]   _zz_5253;
  wire       [15:0]   _zz_5254;
  wire       [15:0]   _zz_5255;
  wire       [15:0]   _zz_5256;
  wire       [15:0]   _zz_5257;
  wire       [15:0]   _zz_5258;
  wire       [15:0]   _zz_5259;
  wire       [15:0]   _zz_5260;
  wire       [15:0]   _zz_5261;
  wire       [15:0]   _zz_5262;
  wire       [15:0]   _zz_5263;
  wire       [15:0]   _zz_5264;
  wire       [31:0]   _zz_5265;
  wire       [31:0]   _zz_5266;
  wire       [15:0]   _zz_5267;
  wire       [31:0]   _zz_5268;
  wire       [31:0]   _zz_5269;
  wire       [15:0]   _zz_5270;
  wire       [15:0]   _zz_5271;
  wire       [15:0]   _zz_5272;
  wire       [15:0]   _zz_5273;
  wire       [15:0]   _zz_5274;
  wire       [15:0]   _zz_5275;
  wire       [15:0]   _zz_5276;
  wire       [15:0]   _zz_5277;
  wire       [15:0]   _zz_5278;
  wire       [15:0]   _zz_5279;
  wire       [15:0]   _zz_5280;
  wire       [15:0]   _zz_5281;
  wire       [15:0]   _zz_5282;
  wire       [15:0]   _zz_5283;
  wire       [15:0]   _zz_5284;
  wire       [15:0]   _zz_5285;
  wire       [15:0]   _zz_5286;
  wire       [31:0]   _zz_5287;
  wire       [31:0]   _zz_5288;
  wire       [15:0]   _zz_5289;
  wire       [31:0]   _zz_5290;
  wire       [31:0]   _zz_5291;
  wire       [15:0]   _zz_5292;
  wire       [15:0]   _zz_5293;
  wire       [15:0]   _zz_5294;
  wire       [15:0]   _zz_5295;
  wire       [15:0]   _zz_5296;
  wire       [15:0]   _zz_5297;
  wire       [15:0]   _zz_5298;
  wire       [15:0]   _zz_5299;
  wire       [15:0]   _zz_5300;
  wire       [15:0]   _zz_5301;
  wire       [15:0]   _zz_5302;
  wire       [15:0]   _zz_5303;
  wire       [15:0]   _zz_5304;
  wire       [15:0]   _zz_5305;
  wire       [15:0]   _zz_5306;
  wire       [15:0]   _zz_5307;
  wire       [15:0]   _zz_5308;
  wire       [31:0]   _zz_5309;
  wire       [31:0]   _zz_5310;
  wire       [15:0]   _zz_5311;
  wire       [31:0]   _zz_5312;
  wire       [31:0]   _zz_5313;
  wire       [15:0]   _zz_5314;
  wire       [15:0]   _zz_5315;
  wire       [15:0]   _zz_5316;
  wire       [15:0]   _zz_5317;
  wire       [15:0]   _zz_5318;
  wire       [15:0]   _zz_5319;
  wire       [15:0]   _zz_5320;
  wire       [15:0]   _zz_5321;
  wire       [15:0]   _zz_5322;
  wire       [15:0]   _zz_5323;
  wire       [15:0]   _zz_5324;
  wire       [15:0]   _zz_5325;
  wire       [15:0]   _zz_5326;
  wire       [15:0]   _zz_5327;
  wire       [15:0]   _zz_5328;
  wire       [15:0]   _zz_5329;
  wire       [15:0]   _zz_5330;
  wire       [31:0]   _zz_5331;
  wire       [31:0]   _zz_5332;
  wire       [15:0]   _zz_5333;
  wire       [31:0]   _zz_5334;
  wire       [31:0]   _zz_5335;
  wire       [15:0]   _zz_5336;
  wire       [15:0]   _zz_5337;
  wire       [15:0]   _zz_5338;
  wire       [15:0]   _zz_5339;
  wire       [15:0]   _zz_5340;
  wire       [15:0]   _zz_5341;
  wire       [15:0]   _zz_5342;
  wire       [15:0]   _zz_5343;
  wire       [15:0]   _zz_5344;
  wire       [15:0]   _zz_5345;
  wire       [15:0]   _zz_5346;
  wire       [15:0]   _zz_5347;
  wire       [15:0]   _zz_5348;
  wire       [15:0]   _zz_5349;
  wire       [15:0]   _zz_5350;
  wire       [15:0]   _zz_5351;
  wire       [15:0]   _zz_5352;
  wire       [31:0]   _zz_5353;
  wire       [31:0]   _zz_5354;
  wire       [15:0]   _zz_5355;
  wire       [31:0]   _zz_5356;
  wire       [31:0]   _zz_5357;
  wire       [15:0]   _zz_5358;
  wire       [15:0]   _zz_5359;
  wire       [15:0]   _zz_5360;
  wire       [15:0]   _zz_5361;
  wire       [15:0]   _zz_5362;
  wire       [15:0]   _zz_5363;
  wire       [15:0]   _zz_5364;
  wire       [15:0]   _zz_5365;
  wire       [15:0]   _zz_5366;
  wire       [15:0]   _zz_5367;
  wire       [15:0]   _zz_5368;
  wire       [15:0]   _zz_5369;
  wire       [15:0]   _zz_5370;
  wire       [15:0]   _zz_5371;
  wire       [15:0]   _zz_5372;
  wire       [15:0]   _zz_5373;
  wire       [15:0]   _zz_5374;
  wire       [31:0]   _zz_5375;
  wire       [31:0]   _zz_5376;
  wire       [15:0]   _zz_5377;
  wire       [31:0]   _zz_5378;
  wire       [31:0]   _zz_5379;
  wire       [15:0]   _zz_5380;
  wire       [15:0]   _zz_5381;
  wire       [15:0]   _zz_5382;
  wire       [15:0]   _zz_5383;
  wire       [15:0]   _zz_5384;
  wire       [15:0]   _zz_5385;
  wire       [15:0]   _zz_5386;
  wire       [15:0]   _zz_5387;
  wire       [15:0]   _zz_5388;
  wire       [15:0]   _zz_5389;
  wire       [15:0]   _zz_5390;
  wire       [15:0]   _zz_5391;
  wire       [15:0]   _zz_5392;
  wire       [15:0]   _zz_5393;
  wire       [15:0]   _zz_5394;
  wire       [15:0]   _zz_5395;
  wire       [15:0]   _zz_5396;
  wire       [31:0]   _zz_5397;
  wire       [31:0]   _zz_5398;
  wire       [15:0]   _zz_5399;
  wire       [31:0]   _zz_5400;
  wire       [31:0]   _zz_5401;
  wire       [15:0]   _zz_5402;
  wire       [15:0]   _zz_5403;
  wire       [15:0]   _zz_5404;
  wire       [15:0]   _zz_5405;
  wire       [15:0]   _zz_5406;
  wire       [15:0]   _zz_5407;
  wire       [15:0]   _zz_5408;
  wire       [15:0]   _zz_5409;
  wire       [15:0]   _zz_5410;
  wire       [15:0]   _zz_5411;
  wire       [15:0]   _zz_5412;
  wire       [15:0]   _zz_5413;
  wire       [15:0]   _zz_5414;
  wire       [15:0]   _zz_5415;
  wire       [15:0]   _zz_5416;
  wire       [15:0]   _zz_5417;
  wire       [15:0]   _zz_5418;
  wire       [31:0]   _zz_5419;
  wire       [31:0]   _zz_5420;
  wire       [15:0]   _zz_5421;
  wire       [31:0]   _zz_5422;
  wire       [31:0]   _zz_5423;
  wire       [15:0]   _zz_5424;
  wire       [15:0]   _zz_5425;
  wire       [15:0]   _zz_5426;
  wire       [15:0]   _zz_5427;
  wire       [15:0]   _zz_5428;
  wire       [15:0]   _zz_5429;
  wire       [15:0]   _zz_5430;
  wire       [15:0]   _zz_5431;
  wire       [15:0]   _zz_5432;
  wire       [15:0]   _zz_5433;
  wire       [15:0]   _zz_5434;
  wire       [15:0]   _zz_5435;
  wire       [15:0]   _zz_5436;
  wire       [15:0]   _zz_5437;
  wire       [15:0]   _zz_5438;
  wire       [15:0]   _zz_5439;
  wire       [15:0]   _zz_5440;
  wire       [31:0]   _zz_5441;
  wire       [31:0]   _zz_5442;
  wire       [15:0]   _zz_5443;
  wire       [31:0]   _zz_5444;
  wire       [31:0]   _zz_5445;
  wire       [15:0]   _zz_5446;
  wire       [15:0]   _zz_5447;
  wire       [15:0]   _zz_5448;
  wire       [15:0]   _zz_5449;
  wire       [15:0]   _zz_5450;
  wire       [15:0]   _zz_5451;
  wire       [15:0]   _zz_5452;
  wire       [15:0]   _zz_5453;
  wire       [15:0]   _zz_5454;
  wire       [15:0]   _zz_5455;
  wire       [15:0]   _zz_5456;
  wire       [15:0]   _zz_5457;
  wire       [15:0]   _zz_5458;
  wire       [15:0]   _zz_5459;
  wire       [15:0]   _zz_5460;
  wire       [15:0]   _zz_5461;
  wire       [15:0]   _zz_5462;
  wire       [31:0]   _zz_5463;
  wire       [31:0]   _zz_5464;
  wire       [15:0]   _zz_5465;
  wire       [31:0]   _zz_5466;
  wire       [31:0]   _zz_5467;
  wire       [15:0]   _zz_5468;
  wire       [15:0]   _zz_5469;
  wire       [15:0]   _zz_5470;
  wire       [15:0]   _zz_5471;
  wire       [15:0]   _zz_5472;
  wire       [15:0]   _zz_5473;
  wire       [15:0]   _zz_5474;
  wire       [15:0]   _zz_5475;
  wire       [15:0]   _zz_5476;
  wire       [15:0]   _zz_5477;
  wire       [15:0]   _zz_5478;
  wire       [15:0]   _zz_5479;
  wire       [15:0]   _zz_5480;
  wire       [15:0]   _zz_5481;
  wire       [15:0]   _zz_5482;
  wire       [15:0]   _zz_5483;
  wire       [15:0]   _zz_5484;
  wire       [31:0]   _zz_5485;
  wire       [31:0]   _zz_5486;
  wire       [15:0]   _zz_5487;
  wire       [31:0]   _zz_5488;
  wire       [31:0]   _zz_5489;
  wire       [15:0]   _zz_5490;
  wire       [15:0]   _zz_5491;
  wire       [15:0]   _zz_5492;
  wire       [15:0]   _zz_5493;
  wire       [15:0]   _zz_5494;
  wire       [15:0]   _zz_5495;
  wire       [15:0]   _zz_5496;
  wire       [15:0]   _zz_5497;
  wire       [15:0]   _zz_5498;
  wire       [15:0]   _zz_5499;
  wire       [15:0]   _zz_5500;
  wire       [15:0]   _zz_5501;
  wire       [15:0]   _zz_5502;
  wire       [15:0]   _zz_5503;
  wire       [15:0]   _zz_5504;
  wire       [15:0]   _zz_5505;
  wire       [15:0]   _zz_5506;
  wire       [31:0]   _zz_5507;
  wire       [31:0]   _zz_5508;
  wire       [15:0]   _zz_5509;
  wire       [31:0]   _zz_5510;
  wire       [31:0]   _zz_5511;
  wire       [15:0]   _zz_5512;
  wire       [15:0]   _zz_5513;
  wire       [15:0]   _zz_5514;
  wire       [15:0]   _zz_5515;
  wire       [15:0]   _zz_5516;
  wire       [15:0]   _zz_5517;
  wire       [15:0]   _zz_5518;
  wire       [15:0]   _zz_5519;
  wire       [15:0]   _zz_5520;
  wire       [15:0]   _zz_5521;
  wire       [15:0]   _zz_5522;
  wire       [15:0]   _zz_5523;
  wire       [15:0]   _zz_5524;
  wire       [15:0]   _zz_5525;
  wire       [15:0]   _zz_5526;
  wire       [15:0]   _zz_5527;
  wire       [15:0]   _zz_5528;
  wire       [31:0]   _zz_5529;
  wire       [31:0]   _zz_5530;
  wire       [15:0]   _zz_5531;
  wire       [31:0]   _zz_5532;
  wire       [31:0]   _zz_5533;
  wire       [15:0]   _zz_5534;
  wire       [15:0]   _zz_5535;
  wire       [15:0]   _zz_5536;
  wire       [15:0]   _zz_5537;
  wire       [15:0]   _zz_5538;
  wire       [15:0]   _zz_5539;
  wire       [15:0]   _zz_5540;
  wire       [15:0]   _zz_5541;
  wire       [15:0]   _zz_5542;
  wire       [15:0]   _zz_5543;
  wire       [15:0]   _zz_5544;
  wire       [15:0]   _zz_5545;
  wire       [15:0]   _zz_5546;
  wire       [15:0]   _zz_5547;
  wire       [15:0]   _zz_5548;
  wire       [15:0]   _zz_5549;
  wire       [15:0]   _zz_5550;
  wire       [31:0]   _zz_5551;
  wire       [31:0]   _zz_5552;
  wire       [15:0]   _zz_5553;
  wire       [31:0]   _zz_5554;
  wire       [31:0]   _zz_5555;
  wire       [15:0]   _zz_5556;
  wire       [15:0]   _zz_5557;
  wire       [15:0]   _zz_5558;
  wire       [15:0]   _zz_5559;
  wire       [15:0]   _zz_5560;
  wire       [15:0]   _zz_5561;
  wire       [15:0]   _zz_5562;
  wire       [15:0]   _zz_5563;
  wire       [15:0]   _zz_5564;
  wire       [15:0]   _zz_5565;
  wire       [15:0]   _zz_5566;
  wire       [15:0]   _zz_5567;
  wire       [15:0]   _zz_5568;
  wire       [15:0]   _zz_5569;
  wire       [15:0]   _zz_5570;
  wire       [15:0]   _zz_5571;
  wire       [15:0]   _zz_5572;
  wire       [31:0]   _zz_5573;
  wire       [31:0]   _zz_5574;
  wire       [15:0]   _zz_5575;
  wire       [31:0]   _zz_5576;
  wire       [31:0]   _zz_5577;
  wire       [15:0]   _zz_5578;
  wire       [15:0]   _zz_5579;
  wire       [15:0]   _zz_5580;
  wire       [15:0]   _zz_5581;
  wire       [15:0]   _zz_5582;
  wire       [15:0]   _zz_5583;
  wire       [15:0]   _zz_5584;
  wire       [15:0]   _zz_5585;
  wire       [15:0]   _zz_5586;
  wire       [15:0]   _zz_5587;
  wire       [15:0]   _zz_5588;
  wire       [15:0]   _zz_5589;
  wire       [15:0]   _zz_5590;
  wire       [15:0]   _zz_5591;
  wire       [15:0]   _zz_5592;
  wire       [15:0]   _zz_5593;
  wire       [15:0]   _zz_5594;
  wire       [31:0]   _zz_5595;
  wire       [31:0]   _zz_5596;
  wire       [15:0]   _zz_5597;
  wire       [31:0]   _zz_5598;
  wire       [31:0]   _zz_5599;
  wire       [15:0]   _zz_5600;
  wire       [15:0]   _zz_5601;
  wire       [15:0]   _zz_5602;
  wire       [15:0]   _zz_5603;
  wire       [15:0]   _zz_5604;
  wire       [15:0]   _zz_5605;
  wire       [15:0]   _zz_5606;
  wire       [15:0]   _zz_5607;
  wire       [15:0]   _zz_5608;
  wire       [15:0]   _zz_5609;
  wire       [15:0]   _zz_5610;
  wire       [15:0]   _zz_5611;
  wire       [15:0]   _zz_5612;
  wire       [15:0]   _zz_5613;
  wire       [15:0]   _zz_5614;
  wire       [15:0]   _zz_5615;
  wire       [15:0]   _zz_5616;
  wire       [31:0]   _zz_5617;
  wire       [31:0]   _zz_5618;
  wire       [15:0]   _zz_5619;
  wire       [31:0]   _zz_5620;
  wire       [31:0]   _zz_5621;
  wire       [15:0]   _zz_5622;
  wire       [15:0]   _zz_5623;
  wire       [15:0]   _zz_5624;
  wire       [15:0]   _zz_5625;
  wire       [15:0]   _zz_5626;
  wire       [15:0]   _zz_5627;
  wire       [15:0]   _zz_5628;
  wire       [15:0]   _zz_5629;
  wire       [15:0]   _zz_5630;
  wire       [15:0]   _zz_5631;
  wire       [15:0]   _zz_5632;
  wire       [15:0]   _zz_5633;
  wire       [15:0]   _zz_5634;
  wire       [15:0]   _zz_5635;
  wire       [15:0]   _zz_5636;
  wire       [15:0]   _zz_5637;
  wire       [15:0]   _zz_5638;
  wire       [31:0]   _zz_5639;
  wire       [31:0]   _zz_5640;
  wire       [15:0]   _zz_5641;
  wire       [31:0]   _zz_5642;
  wire       [31:0]   _zz_5643;
  wire       [15:0]   _zz_5644;
  wire       [15:0]   _zz_5645;
  wire       [15:0]   _zz_5646;
  wire       [15:0]   _zz_5647;
  wire       [15:0]   _zz_5648;
  wire       [15:0]   _zz_5649;
  wire       [15:0]   _zz_5650;
  wire       [15:0]   _zz_5651;
  wire       [15:0]   _zz_5652;
  wire       [15:0]   _zz_5653;
  wire       [15:0]   _zz_5654;
  wire       [15:0]   _zz_5655;
  wire       [15:0]   _zz_5656;
  wire       [15:0]   _zz_5657;
  wire       [15:0]   _zz_5658;
  wire       [15:0]   _zz_5659;
  wire       [15:0]   _zz_5660;
  wire       [31:0]   _zz_5661;
  wire       [31:0]   _zz_5662;
  wire       [15:0]   _zz_5663;
  wire       [31:0]   _zz_5664;
  wire       [31:0]   _zz_5665;
  wire       [15:0]   _zz_5666;
  wire       [15:0]   _zz_5667;
  wire       [15:0]   _zz_5668;
  wire       [15:0]   _zz_5669;
  wire       [15:0]   _zz_5670;
  wire       [15:0]   _zz_5671;
  wire       [15:0]   _zz_5672;
  wire       [15:0]   _zz_5673;
  wire       [15:0]   _zz_5674;
  wire       [15:0]   _zz_5675;
  wire       [15:0]   _zz_5676;
  wire       [15:0]   _zz_5677;
  wire       [15:0]   _zz_5678;
  wire       [15:0]   _zz_5679;
  wire       [15:0]   _zz_5680;
  wire       [15:0]   _zz_5681;
  wire       [15:0]   _zz_5682;
  wire       [31:0]   _zz_5683;
  wire       [31:0]   _zz_5684;
  wire       [15:0]   _zz_5685;
  wire       [31:0]   _zz_5686;
  wire       [31:0]   _zz_5687;
  wire       [15:0]   _zz_5688;
  wire       [15:0]   _zz_5689;
  wire       [15:0]   _zz_5690;
  wire       [15:0]   _zz_5691;
  wire       [15:0]   _zz_5692;
  wire       [15:0]   _zz_5693;
  wire       [15:0]   _zz_5694;
  wire       [15:0]   _zz_5695;
  wire       [15:0]   _zz_5696;
  wire       [15:0]   _zz_5697;
  wire       [15:0]   _zz_5698;
  wire       [15:0]   _zz_5699;
  wire       [15:0]   _zz_5700;
  wire       [15:0]   _zz_5701;
  wire       [15:0]   _zz_5702;
  wire       [15:0]   _zz_5703;
  wire       [15:0]   _zz_5704;
  wire       [31:0]   _zz_5705;
  wire       [31:0]   _zz_5706;
  wire       [15:0]   _zz_5707;
  wire       [31:0]   _zz_5708;
  wire       [31:0]   _zz_5709;
  wire       [15:0]   _zz_5710;
  wire       [15:0]   _zz_5711;
  wire       [15:0]   _zz_5712;
  wire       [15:0]   _zz_5713;
  wire       [15:0]   _zz_5714;
  wire       [15:0]   _zz_5715;
  wire       [15:0]   _zz_5716;
  wire       [15:0]   _zz_5717;
  wire       [15:0]   _zz_5718;
  wire       [15:0]   _zz_5719;
  wire       [15:0]   _zz_5720;
  wire       [15:0]   _zz_5721;
  wire       [15:0]   _zz_5722;
  wire       [15:0]   _zz_5723;
  wire       [15:0]   _zz_5724;
  wire       [15:0]   _zz_5725;
  wire       [15:0]   _zz_5726;
  wire       [31:0]   _zz_5727;
  wire       [31:0]   _zz_5728;
  wire       [15:0]   _zz_5729;
  wire       [31:0]   _zz_5730;
  wire       [31:0]   _zz_5731;
  wire       [15:0]   _zz_5732;
  wire       [15:0]   _zz_5733;
  wire       [15:0]   _zz_5734;
  wire       [15:0]   _zz_5735;
  wire       [15:0]   _zz_5736;
  wire       [15:0]   _zz_5737;
  wire       [15:0]   _zz_5738;
  wire       [15:0]   _zz_5739;
  wire       [15:0]   _zz_5740;
  wire       [15:0]   _zz_5741;
  wire       [15:0]   _zz_5742;
  wire       [15:0]   _zz_5743;
  wire       [15:0]   _zz_5744;
  wire       [15:0]   _zz_5745;
  wire       [15:0]   _zz_5746;
  wire       [15:0]   _zz_5747;
  wire       [15:0]   _zz_5748;
  wire       [31:0]   _zz_5749;
  wire       [31:0]   _zz_5750;
  wire       [15:0]   _zz_5751;
  wire       [31:0]   _zz_5752;
  wire       [31:0]   _zz_5753;
  wire       [15:0]   _zz_5754;
  wire       [15:0]   _zz_5755;
  wire       [15:0]   _zz_5756;
  wire       [15:0]   _zz_5757;
  wire       [15:0]   _zz_5758;
  wire       [15:0]   _zz_5759;
  wire       [15:0]   _zz_5760;
  wire       [15:0]   _zz_5761;
  wire       [15:0]   _zz_5762;
  wire       [15:0]   _zz_5763;
  wire       [15:0]   _zz_5764;
  wire       [15:0]   _zz_5765;
  wire       [15:0]   _zz_5766;
  wire       [15:0]   _zz_5767;
  wire       [15:0]   _zz_5768;
  wire       [15:0]   _zz_5769;
  wire       [15:0]   _zz_5770;
  wire       [31:0]   _zz_5771;
  wire       [31:0]   _zz_5772;
  wire       [15:0]   _zz_5773;
  wire       [31:0]   _zz_5774;
  wire       [31:0]   _zz_5775;
  wire       [15:0]   _zz_5776;
  wire       [15:0]   _zz_5777;
  wire       [15:0]   _zz_5778;
  wire       [15:0]   _zz_5779;
  wire       [15:0]   _zz_5780;
  wire       [15:0]   _zz_5781;
  wire       [15:0]   _zz_5782;
  wire       [15:0]   _zz_5783;
  wire       [15:0]   _zz_5784;
  wire       [15:0]   _zz_5785;
  wire       [15:0]   _zz_5786;
  wire       [15:0]   _zz_5787;
  wire       [15:0]   _zz_5788;
  wire       [15:0]   _zz_5789;
  wire       [15:0]   _zz_5790;
  wire       [15:0]   _zz_5791;
  wire       [15:0]   _zz_5792;
  wire       [31:0]   _zz_5793;
  wire       [31:0]   _zz_5794;
  wire       [15:0]   _zz_5795;
  wire       [31:0]   _zz_5796;
  wire       [31:0]   _zz_5797;
  wire       [15:0]   _zz_5798;
  wire       [15:0]   _zz_5799;
  wire       [15:0]   _zz_5800;
  wire       [15:0]   _zz_5801;
  wire       [15:0]   _zz_5802;
  wire       [15:0]   _zz_5803;
  wire       [15:0]   _zz_5804;
  wire       [15:0]   _zz_5805;
  wire       [15:0]   _zz_5806;
  wire       [15:0]   _zz_5807;
  wire       [15:0]   _zz_5808;
  wire       [15:0]   _zz_5809;
  wire       [15:0]   _zz_5810;
  wire       [15:0]   _zz_5811;
  wire       [15:0]   _zz_5812;
  wire       [15:0]   _zz_5813;
  wire       [15:0]   _zz_5814;
  wire       [31:0]   _zz_5815;
  wire       [31:0]   _zz_5816;
  wire       [15:0]   _zz_5817;
  wire       [31:0]   _zz_5818;
  wire       [31:0]   _zz_5819;
  wire       [15:0]   _zz_5820;
  wire       [15:0]   _zz_5821;
  wire       [15:0]   _zz_5822;
  wire       [15:0]   _zz_5823;
  wire       [15:0]   _zz_5824;
  wire       [15:0]   _zz_5825;
  wire       [15:0]   _zz_5826;
  wire       [15:0]   _zz_5827;
  wire       [15:0]   _zz_5828;
  wire       [15:0]   _zz_5829;
  wire       [15:0]   _zz_5830;
  wire       [15:0]   _zz_5831;
  wire       [15:0]   _zz_5832;
  wire       [15:0]   _zz_5833;
  wire       [15:0]   _zz_5834;
  wire       [15:0]   _zz_5835;
  wire       [15:0]   _zz_5836;
  wire       [31:0]   _zz_5837;
  wire       [31:0]   _zz_5838;
  wire       [15:0]   _zz_5839;
  wire       [31:0]   _zz_5840;
  wire       [31:0]   _zz_5841;
  wire       [15:0]   _zz_5842;
  wire       [15:0]   _zz_5843;
  wire       [15:0]   _zz_5844;
  wire       [15:0]   _zz_5845;
  wire       [15:0]   _zz_5846;
  wire       [15:0]   _zz_5847;
  wire       [15:0]   _zz_5848;
  wire       [15:0]   _zz_5849;
  wire       [15:0]   _zz_5850;
  wire       [15:0]   _zz_5851;
  wire       [15:0]   _zz_5852;
  wire       [15:0]   _zz_5853;
  wire       [15:0]   _zz_5854;
  wire       [15:0]   _zz_5855;
  wire       [15:0]   _zz_5856;
  wire       [15:0]   _zz_5857;
  wire       [15:0]   _zz_5858;
  wire       [31:0]   _zz_5859;
  wire       [31:0]   _zz_5860;
  wire       [15:0]   _zz_5861;
  wire       [31:0]   _zz_5862;
  wire       [31:0]   _zz_5863;
  wire       [15:0]   _zz_5864;
  wire       [15:0]   _zz_5865;
  wire       [15:0]   _zz_5866;
  wire       [15:0]   _zz_5867;
  wire       [15:0]   _zz_5868;
  wire       [15:0]   _zz_5869;
  wire       [15:0]   _zz_5870;
  wire       [15:0]   _zz_5871;
  wire       [15:0]   _zz_5872;
  wire       [15:0]   _zz_5873;
  wire       [15:0]   _zz_5874;
  wire       [15:0]   _zz_5875;
  wire       [15:0]   _zz_5876;
  wire       [15:0]   _zz_5877;
  wire       [15:0]   _zz_5878;
  wire       [15:0]   _zz_5879;
  wire       [15:0]   _zz_5880;
  wire       [31:0]   _zz_5881;
  wire       [31:0]   _zz_5882;
  wire       [15:0]   _zz_5883;
  wire       [31:0]   _zz_5884;
  wire       [31:0]   _zz_5885;
  wire       [15:0]   _zz_5886;
  wire       [15:0]   _zz_5887;
  wire       [15:0]   _zz_5888;
  wire       [15:0]   _zz_5889;
  wire       [15:0]   _zz_5890;
  wire       [15:0]   _zz_5891;
  wire       [15:0]   _zz_5892;
  wire       [15:0]   _zz_5893;
  wire       [15:0]   _zz_5894;
  wire       [15:0]   _zz_5895;
  wire       [15:0]   _zz_5896;
  wire       [15:0]   _zz_5897;
  wire       [15:0]   _zz_5898;
  wire       [15:0]   _zz_5899;
  wire       [15:0]   _zz_5900;
  wire       [15:0]   _zz_5901;
  wire       [15:0]   _zz_5902;
  wire       [31:0]   _zz_5903;
  wire       [31:0]   _zz_5904;
  wire       [15:0]   _zz_5905;
  wire       [31:0]   _zz_5906;
  wire       [31:0]   _zz_5907;
  wire       [15:0]   _zz_5908;
  wire       [15:0]   _zz_5909;
  wire       [15:0]   _zz_5910;
  wire       [15:0]   _zz_5911;
  wire       [15:0]   _zz_5912;
  wire       [15:0]   _zz_5913;
  wire       [15:0]   _zz_5914;
  wire       [15:0]   _zz_5915;
  wire       [15:0]   _zz_5916;
  wire       [15:0]   _zz_5917;
  wire       [15:0]   _zz_5918;
  wire       [15:0]   _zz_5919;
  wire       [15:0]   _zz_5920;
  wire       [15:0]   _zz_5921;
  wire       [15:0]   _zz_5922;
  wire       [15:0]   _zz_5923;
  wire       [15:0]   _zz_5924;
  wire       [31:0]   _zz_5925;
  wire       [31:0]   _zz_5926;
  wire       [15:0]   _zz_5927;
  wire       [31:0]   _zz_5928;
  wire       [31:0]   _zz_5929;
  wire       [15:0]   _zz_5930;
  wire       [15:0]   _zz_5931;
  wire       [15:0]   _zz_5932;
  wire       [15:0]   _zz_5933;
  wire       [15:0]   _zz_5934;
  wire       [15:0]   _zz_5935;
  wire       [15:0]   _zz_5936;
  wire       [15:0]   _zz_5937;
  wire       [15:0]   _zz_5938;
  wire       [15:0]   _zz_5939;
  wire       [15:0]   _zz_5940;
  wire       [15:0]   _zz_5941;
  wire       [15:0]   _zz_5942;
  wire       [15:0]   _zz_5943;
  wire       [15:0]   _zz_5944;
  wire       [15:0]   _zz_5945;
  wire       [15:0]   _zz_5946;
  wire       [31:0]   _zz_5947;
  wire       [31:0]   _zz_5948;
  wire       [15:0]   _zz_5949;
  wire       [31:0]   _zz_5950;
  wire       [31:0]   _zz_5951;
  wire       [15:0]   _zz_5952;
  wire       [15:0]   _zz_5953;
  wire       [15:0]   _zz_5954;
  wire       [15:0]   _zz_5955;
  wire       [15:0]   _zz_5956;
  wire       [15:0]   _zz_5957;
  wire       [15:0]   _zz_5958;
  wire       [15:0]   _zz_5959;
  wire       [15:0]   _zz_5960;
  wire       [15:0]   _zz_5961;
  wire       [15:0]   _zz_5962;
  wire       [15:0]   _zz_5963;
  wire       [15:0]   _zz_5964;
  wire       [15:0]   _zz_5965;
  wire       [15:0]   _zz_5966;
  wire       [15:0]   _zz_5967;
  wire       [15:0]   _zz_5968;
  wire       [31:0]   _zz_5969;
  wire       [31:0]   _zz_5970;
  wire       [15:0]   _zz_5971;
  wire       [31:0]   _zz_5972;
  wire       [31:0]   _zz_5973;
  wire       [15:0]   _zz_5974;
  wire       [15:0]   _zz_5975;
  wire       [15:0]   _zz_5976;
  wire       [15:0]   _zz_5977;
  wire       [15:0]   _zz_5978;
  wire       [15:0]   _zz_5979;
  wire       [15:0]   _zz_5980;
  wire       [15:0]   _zz_5981;
  wire       [15:0]   _zz_5982;
  wire       [15:0]   _zz_5983;
  wire       [15:0]   _zz_5984;
  wire       [15:0]   _zz_5985;
  wire       [15:0]   _zz_5986;
  wire       [15:0]   _zz_5987;
  wire       [15:0]   _zz_5988;
  wire       [15:0]   _zz_5989;
  wire       [15:0]   _zz_5990;
  wire       [31:0]   _zz_5991;
  wire       [31:0]   _zz_5992;
  wire       [15:0]   _zz_5993;
  wire       [31:0]   _zz_5994;
  wire       [31:0]   _zz_5995;
  wire       [15:0]   _zz_5996;
  wire       [15:0]   _zz_5997;
  wire       [15:0]   _zz_5998;
  wire       [15:0]   _zz_5999;
  wire       [15:0]   _zz_6000;
  wire       [15:0]   _zz_6001;
  wire       [15:0]   _zz_6002;
  wire       [15:0]   _zz_6003;
  wire       [15:0]   _zz_6004;
  wire       [15:0]   _zz_6005;
  wire       [15:0]   _zz_6006;
  wire       [15:0]   _zz_6007;
  wire       [15:0]   _zz_6008;
  wire       [15:0]   _zz_6009;
  wire       [15:0]   _zz_6010;
  wire       [15:0]   _zz_6011;
  wire       [15:0]   _zz_6012;
  wire       [31:0]   _zz_6013;
  wire       [31:0]   _zz_6014;
  wire       [15:0]   _zz_6015;
  wire       [31:0]   _zz_6016;
  wire       [31:0]   _zz_6017;
  wire       [15:0]   _zz_6018;
  wire       [15:0]   _zz_6019;
  wire       [15:0]   _zz_6020;
  wire       [15:0]   _zz_6021;
  wire       [15:0]   _zz_6022;
  wire       [15:0]   _zz_6023;
  wire       [15:0]   _zz_6024;
  wire       [15:0]   _zz_6025;
  wire       [15:0]   _zz_6026;
  wire       [15:0]   _zz_6027;
  wire       [15:0]   _zz_6028;
  wire       [15:0]   _zz_6029;
  wire       [15:0]   _zz_6030;
  wire       [15:0]   _zz_6031;
  wire       [15:0]   _zz_6032;
  wire       [15:0]   _zz_6033;
  wire       [15:0]   _zz_6034;
  wire       [31:0]   _zz_6035;
  wire       [31:0]   _zz_6036;
  wire       [15:0]   _zz_6037;
  wire       [31:0]   _zz_6038;
  wire       [31:0]   _zz_6039;
  wire       [15:0]   _zz_6040;
  wire       [15:0]   _zz_6041;
  wire       [15:0]   _zz_6042;
  wire       [15:0]   _zz_6043;
  wire       [15:0]   _zz_6044;
  wire       [15:0]   _zz_6045;
  wire       [15:0]   _zz_6046;
  wire       [15:0]   _zz_6047;
  wire       [15:0]   _zz_6048;
  wire       [15:0]   _zz_6049;
  wire       [15:0]   _zz_6050;
  wire       [15:0]   _zz_6051;
  wire       [15:0]   _zz_6052;
  wire       [15:0]   _zz_6053;
  wire       [15:0]   _zz_6054;
  wire       [15:0]   _zz_6055;
  wire       [15:0]   _zz_6056;
  wire       [31:0]   _zz_6057;
  wire       [31:0]   _zz_6058;
  wire       [15:0]   _zz_6059;
  wire       [31:0]   _zz_6060;
  wire       [31:0]   _zz_6061;
  wire       [15:0]   _zz_6062;
  wire       [15:0]   _zz_6063;
  wire       [15:0]   _zz_6064;
  wire       [15:0]   _zz_6065;
  wire       [15:0]   _zz_6066;
  wire       [15:0]   _zz_6067;
  wire       [15:0]   _zz_6068;
  wire       [15:0]   _zz_6069;
  wire       [15:0]   _zz_6070;
  wire       [15:0]   _zz_6071;
  wire       [15:0]   _zz_6072;
  wire       [15:0]   _zz_6073;
  wire       [15:0]   _zz_6074;
  wire       [15:0]   _zz_6075;
  wire       [15:0]   _zz_6076;
  wire       [15:0]   _zz_6077;
  wire       [15:0]   _zz_6078;
  wire       [31:0]   _zz_6079;
  wire       [31:0]   _zz_6080;
  wire       [15:0]   _zz_6081;
  wire       [31:0]   _zz_6082;
  wire       [31:0]   _zz_6083;
  wire       [15:0]   _zz_6084;
  wire       [15:0]   _zz_6085;
  wire       [15:0]   _zz_6086;
  wire       [15:0]   _zz_6087;
  wire       [15:0]   _zz_6088;
  wire       [15:0]   _zz_6089;
  wire       [15:0]   _zz_6090;
  wire       [15:0]   _zz_6091;
  wire       [15:0]   _zz_6092;
  wire       [15:0]   _zz_6093;
  wire       [15:0]   _zz_6094;
  wire       [15:0]   _zz_6095;
  wire       [15:0]   _zz_6096;
  wire       [15:0]   _zz_6097;
  wire       [15:0]   _zz_6098;
  wire       [15:0]   _zz_6099;
  wire       [15:0]   _zz_6100;
  wire       [31:0]   _zz_6101;
  wire       [31:0]   _zz_6102;
  wire       [15:0]   _zz_6103;
  wire       [31:0]   _zz_6104;
  wire       [31:0]   _zz_6105;
  wire       [15:0]   _zz_6106;
  wire       [15:0]   _zz_6107;
  wire       [15:0]   _zz_6108;
  wire       [15:0]   _zz_6109;
  wire       [15:0]   _zz_6110;
  wire       [15:0]   _zz_6111;
  wire       [15:0]   _zz_6112;
  wire       [15:0]   _zz_6113;
  wire       [15:0]   _zz_6114;
  wire       [15:0]   _zz_6115;
  wire       [15:0]   _zz_6116;
  wire       [15:0]   _zz_6117;
  wire       [15:0]   _zz_6118;
  wire       [15:0]   _zz_6119;
  wire       [15:0]   _zz_6120;
  wire       [15:0]   _zz_6121;
  wire       [15:0]   _zz_6122;
  wire       [31:0]   _zz_6123;
  wire       [31:0]   _zz_6124;
  wire       [15:0]   _zz_6125;
  wire       [31:0]   _zz_6126;
  wire       [31:0]   _zz_6127;
  wire       [15:0]   _zz_6128;
  wire       [15:0]   _zz_6129;
  wire       [15:0]   _zz_6130;
  wire       [15:0]   _zz_6131;
  wire       [15:0]   _zz_6132;
  wire       [15:0]   _zz_6133;
  wire       [15:0]   _zz_6134;
  wire       [15:0]   _zz_6135;
  wire       [15:0]   _zz_6136;
  wire       [15:0]   _zz_6137;
  wire       [15:0]   _zz_6138;
  wire       [15:0]   _zz_6139;
  wire       [15:0]   _zz_6140;
  wire       [15:0]   _zz_6141;
  wire       [15:0]   _zz_6142;
  wire       [15:0]   _zz_6143;
  wire       [15:0]   _zz_6144;
  wire       [31:0]   _zz_6145;
  wire       [31:0]   _zz_6146;
  wire       [15:0]   _zz_6147;
  wire       [31:0]   _zz_6148;
  wire       [31:0]   _zz_6149;
  wire       [15:0]   _zz_6150;
  wire       [15:0]   _zz_6151;
  wire       [15:0]   _zz_6152;
  wire       [15:0]   _zz_6153;
  wire       [15:0]   _zz_6154;
  wire       [15:0]   _zz_6155;
  wire       [15:0]   _zz_6156;
  wire       [15:0]   _zz_6157;
  wire       [15:0]   _zz_6158;
  wire       [15:0]   _zz_6159;
  wire       [15:0]   _zz_6160;
  wire       [15:0]   _zz_6161;
  wire       [15:0]   _zz_6162;
  wire       [15:0]   _zz_6163;
  wire       [15:0]   _zz_6164;
  wire       [15:0]   _zz_6165;
  wire       [15:0]   _zz_6166;
  wire       [31:0]   _zz_6167;
  wire       [31:0]   _zz_6168;
  wire       [15:0]   _zz_6169;
  wire       [31:0]   _zz_6170;
  wire       [31:0]   _zz_6171;
  wire       [15:0]   _zz_6172;
  wire       [15:0]   _zz_6173;
  wire       [15:0]   _zz_6174;
  wire       [15:0]   _zz_6175;
  wire       [15:0]   _zz_6176;
  wire       [15:0]   _zz_6177;
  wire       [15:0]   _zz_6178;
  wire       [15:0]   _zz_6179;
  wire       [15:0]   _zz_6180;
  wire       [15:0]   _zz_6181;
  wire       [15:0]   _zz_6182;
  wire       [15:0]   _zz_6183;
  wire       [15:0]   _zz_6184;
  wire       [15:0]   _zz_6185;
  wire       [15:0]   _zz_6186;
  wire       [15:0]   _zz_6187;
  wire       [15:0]   _zz_6188;
  wire       [31:0]   _zz_6189;
  wire       [31:0]   _zz_6190;
  wire       [15:0]   _zz_6191;
  wire       [31:0]   _zz_6192;
  wire       [31:0]   _zz_6193;
  wire       [15:0]   _zz_6194;
  wire       [15:0]   _zz_6195;
  wire       [15:0]   _zz_6196;
  wire       [15:0]   _zz_6197;
  wire       [15:0]   _zz_6198;
  wire       [15:0]   _zz_6199;
  wire       [15:0]   _zz_6200;
  wire       [15:0]   _zz_6201;
  wire       [15:0]   _zz_6202;
  wire       [15:0]   _zz_6203;
  wire       [15:0]   _zz_6204;
  wire       [15:0]   _zz_6205;
  wire       [15:0]   _zz_6206;
  wire       [15:0]   _zz_6207;
  wire       [15:0]   _zz_6208;
  wire       [15:0]   _zz_6209;
  wire       [15:0]   _zz_6210;
  wire       [31:0]   _zz_6211;
  wire       [31:0]   _zz_6212;
  wire       [15:0]   _zz_6213;
  wire       [31:0]   _zz_6214;
  wire       [31:0]   _zz_6215;
  wire       [15:0]   _zz_6216;
  wire       [15:0]   _zz_6217;
  wire       [15:0]   _zz_6218;
  wire       [15:0]   _zz_6219;
  wire       [15:0]   _zz_6220;
  wire       [15:0]   _zz_6221;
  wire       [15:0]   _zz_6222;
  wire       [15:0]   _zz_6223;
  wire       [15:0]   _zz_6224;
  wire       [15:0]   _zz_6225;
  wire       [15:0]   _zz_6226;
  wire       [15:0]   _zz_6227;
  wire       [15:0]   _zz_6228;
  wire       [15:0]   _zz_6229;
  wire       [15:0]   _zz_6230;
  wire       [15:0]   _zz_6231;
  wire       [15:0]   _zz_6232;
  wire       [31:0]   _zz_6233;
  wire       [31:0]   _zz_6234;
  wire       [15:0]   _zz_6235;
  wire       [31:0]   _zz_6236;
  wire       [31:0]   _zz_6237;
  wire       [15:0]   _zz_6238;
  wire       [15:0]   _zz_6239;
  wire       [15:0]   _zz_6240;
  wire       [15:0]   _zz_6241;
  wire       [15:0]   _zz_6242;
  wire       [15:0]   _zz_6243;
  wire       [15:0]   _zz_6244;
  wire       [15:0]   _zz_6245;
  wire       [15:0]   _zz_6246;
  wire       [15:0]   _zz_6247;
  wire       [15:0]   _zz_6248;
  wire       [15:0]   _zz_6249;
  wire       [15:0]   _zz_6250;
  wire       [15:0]   _zz_6251;
  wire       [15:0]   _zz_6252;
  wire       [15:0]   _zz_6253;
  wire       [15:0]   _zz_6254;
  wire       [31:0]   _zz_6255;
  wire       [31:0]   _zz_6256;
  wire       [15:0]   _zz_6257;
  wire       [31:0]   _zz_6258;
  wire       [31:0]   _zz_6259;
  wire       [15:0]   _zz_6260;
  wire       [15:0]   _zz_6261;
  wire       [15:0]   _zz_6262;
  wire       [15:0]   _zz_6263;
  wire       [15:0]   _zz_6264;
  wire       [15:0]   _zz_6265;
  wire       [15:0]   _zz_6266;
  wire       [15:0]   _zz_6267;
  wire       [15:0]   _zz_6268;
  wire       [15:0]   _zz_6269;
  wire       [15:0]   _zz_6270;
  wire       [15:0]   _zz_6271;
  wire       [15:0]   _zz_6272;
  wire       [15:0]   _zz_6273;
  wire       [15:0]   _zz_6274;
  wire       [15:0]   _zz_6275;
  wire       [15:0]   _zz_6276;
  wire       [31:0]   _zz_6277;
  wire       [31:0]   _zz_6278;
  wire       [15:0]   _zz_6279;
  wire       [31:0]   _zz_6280;
  wire       [31:0]   _zz_6281;
  wire       [15:0]   _zz_6282;
  wire       [15:0]   _zz_6283;
  wire       [15:0]   _zz_6284;
  wire       [15:0]   _zz_6285;
  wire       [15:0]   _zz_6286;
  wire       [15:0]   _zz_6287;
  wire       [15:0]   _zz_6288;
  wire       [15:0]   _zz_6289;
  wire       [15:0]   _zz_6290;
  wire       [15:0]   _zz_6291;
  wire       [15:0]   _zz_6292;
  wire       [15:0]   _zz_6293;
  wire       [15:0]   _zz_6294;
  wire       [15:0]   _zz_6295;
  wire       [15:0]   _zz_6296;
  wire       [15:0]   _zz_6297;
  wire       [15:0]   _zz_6298;
  wire       [31:0]   _zz_6299;
  wire       [31:0]   _zz_6300;
  wire       [15:0]   _zz_6301;
  wire       [31:0]   _zz_6302;
  wire       [31:0]   _zz_6303;
  wire       [15:0]   _zz_6304;
  wire       [15:0]   _zz_6305;
  wire       [15:0]   _zz_6306;
  wire       [15:0]   _zz_6307;
  wire       [15:0]   _zz_6308;
  wire       [15:0]   _zz_6309;
  wire       [15:0]   _zz_6310;
  wire       [15:0]   _zz_6311;
  wire       [15:0]   _zz_6312;
  wire       [15:0]   _zz_6313;
  wire       [15:0]   _zz_6314;
  wire       [15:0]   _zz_6315;
  wire       [15:0]   _zz_6316;
  wire       [15:0]   _zz_6317;
  wire       [15:0]   _zz_6318;
  wire       [15:0]   _zz_6319;
  wire       [15:0]   _zz_6320;
  wire       [31:0]   _zz_6321;
  wire       [31:0]   _zz_6322;
  wire       [15:0]   _zz_6323;
  wire       [31:0]   _zz_6324;
  wire       [31:0]   _zz_6325;
  wire       [15:0]   _zz_6326;
  wire       [15:0]   _zz_6327;
  wire       [15:0]   _zz_6328;
  wire       [15:0]   _zz_6329;
  wire       [15:0]   _zz_6330;
  wire       [15:0]   _zz_6331;
  wire       [15:0]   _zz_6332;
  wire       [15:0]   _zz_6333;
  wire       [15:0]   _zz_6334;
  wire       [15:0]   _zz_6335;
  wire       [15:0]   _zz_6336;
  wire       [15:0]   _zz_6337;
  wire       [15:0]   _zz_6338;
  wire       [15:0]   _zz_6339;
  wire       [15:0]   _zz_6340;
  wire       [15:0]   _zz_6341;
  wire       [15:0]   _zz_6342;
  wire       [31:0]   _zz_6343;
  wire       [31:0]   _zz_6344;
  wire       [15:0]   _zz_6345;
  wire       [31:0]   _zz_6346;
  wire       [31:0]   _zz_6347;
  wire       [15:0]   _zz_6348;
  wire       [15:0]   _zz_6349;
  wire       [15:0]   _zz_6350;
  wire       [15:0]   _zz_6351;
  wire       [15:0]   _zz_6352;
  wire       [15:0]   _zz_6353;
  wire       [15:0]   _zz_6354;
  wire       [15:0]   _zz_6355;
  wire       [15:0]   _zz_6356;
  wire       [15:0]   _zz_6357;
  wire       [15:0]   _zz_6358;
  wire       [15:0]   _zz_6359;
  wire       [15:0]   _zz_6360;
  wire       [15:0]   _zz_6361;
  wire       [15:0]   _zz_6362;
  wire       [15:0]   _zz_6363;
  wire       [15:0]   _zz_6364;
  wire       [31:0]   _zz_6365;
  wire       [31:0]   _zz_6366;
  wire       [15:0]   _zz_6367;
  wire       [31:0]   _zz_6368;
  wire       [31:0]   _zz_6369;
  wire       [15:0]   _zz_6370;
  wire       [15:0]   _zz_6371;
  wire       [15:0]   _zz_6372;
  wire       [15:0]   _zz_6373;
  wire       [15:0]   _zz_6374;
  wire       [15:0]   _zz_6375;
  wire       [15:0]   _zz_6376;
  wire       [15:0]   _zz_6377;
  wire       [15:0]   _zz_6378;
  wire       [15:0]   _zz_6379;
  wire       [15:0]   _zz_6380;
  wire       [15:0]   _zz_6381;
  wire       [15:0]   _zz_6382;
  wire       [15:0]   _zz_6383;
  wire       [15:0]   _zz_6384;
  wire       [15:0]   _zz_6385;
  wire       [15:0]   _zz_6386;
  wire       [31:0]   _zz_6387;
  wire       [31:0]   _zz_6388;
  wire       [15:0]   _zz_6389;
  wire       [31:0]   _zz_6390;
  wire       [31:0]   _zz_6391;
  wire       [15:0]   _zz_6392;
  wire       [15:0]   _zz_6393;
  wire       [15:0]   _zz_6394;
  wire       [15:0]   _zz_6395;
  wire       [15:0]   _zz_6396;
  wire       [15:0]   _zz_6397;
  wire       [15:0]   _zz_6398;
  wire       [15:0]   _zz_6399;
  wire       [15:0]   _zz_6400;
  wire       [15:0]   _zz_6401;
  wire       [15:0]   _zz_6402;
  wire       [15:0]   _zz_6403;
  wire       [15:0]   _zz_6404;
  wire       [15:0]   _zz_6405;
  wire       [15:0]   _zz_6406;
  wire       [15:0]   _zz_6407;
  wire       [15:0]   _zz_6408;
  wire       [31:0]   _zz_6409;
  wire       [31:0]   _zz_6410;
  wire       [15:0]   _zz_6411;
  wire       [31:0]   _zz_6412;
  wire       [31:0]   _zz_6413;
  wire       [15:0]   _zz_6414;
  wire       [15:0]   _zz_6415;
  wire       [15:0]   _zz_6416;
  wire       [15:0]   _zz_6417;
  wire       [15:0]   _zz_6418;
  wire       [15:0]   _zz_6419;
  wire       [15:0]   _zz_6420;
  wire       [15:0]   _zz_6421;
  wire       [15:0]   _zz_6422;
  wire       [15:0]   _zz_6423;
  wire       [15:0]   _zz_6424;
  wire       [15:0]   _zz_6425;
  wire       [15:0]   _zz_6426;
  wire       [15:0]   _zz_6427;
  wire       [15:0]   _zz_6428;
  wire       [15:0]   _zz_6429;
  wire       [15:0]   _zz_6430;
  wire       [31:0]   _zz_6431;
  wire       [31:0]   _zz_6432;
  wire       [15:0]   _zz_6433;
  wire       [31:0]   _zz_6434;
  wire       [31:0]   _zz_6435;
  wire       [15:0]   _zz_6436;
  wire       [15:0]   _zz_6437;
  wire       [15:0]   _zz_6438;
  wire       [15:0]   _zz_6439;
  wire       [15:0]   _zz_6440;
  wire       [15:0]   _zz_6441;
  wire       [15:0]   _zz_6442;
  wire       [15:0]   _zz_6443;
  wire       [15:0]   _zz_6444;
  wire       [15:0]   _zz_6445;
  wire       [15:0]   _zz_6446;
  wire       [15:0]   _zz_6447;
  wire       [15:0]   _zz_6448;
  wire       [15:0]   _zz_6449;
  wire       [15:0]   _zz_6450;
  wire       [15:0]   _zz_6451;
  wire       [15:0]   _zz_6452;
  wire       [31:0]   _zz_6453;
  wire       [31:0]   _zz_6454;
  wire       [15:0]   _zz_6455;
  wire       [31:0]   _zz_6456;
  wire       [31:0]   _zz_6457;
  wire       [15:0]   _zz_6458;
  wire       [15:0]   _zz_6459;
  wire       [15:0]   _zz_6460;
  wire       [15:0]   _zz_6461;
  wire       [15:0]   _zz_6462;
  wire       [15:0]   _zz_6463;
  wire       [15:0]   _zz_6464;
  wire       [15:0]   _zz_6465;
  wire       [15:0]   _zz_6466;
  wire       [15:0]   _zz_6467;
  wire       [15:0]   _zz_6468;
  wire       [15:0]   _zz_6469;
  wire       [15:0]   _zz_6470;
  wire       [15:0]   _zz_6471;
  wire       [15:0]   _zz_6472;
  wire       [15:0]   _zz_6473;
  wire       [15:0]   _zz_6474;
  wire       [31:0]   _zz_6475;
  wire       [31:0]   _zz_6476;
  wire       [15:0]   _zz_6477;
  wire       [31:0]   _zz_6478;
  wire       [31:0]   _zz_6479;
  wire       [15:0]   _zz_6480;
  wire       [15:0]   _zz_6481;
  wire       [15:0]   _zz_6482;
  wire       [15:0]   _zz_6483;
  wire       [15:0]   _zz_6484;
  wire       [15:0]   _zz_6485;
  wire       [15:0]   _zz_6486;
  wire       [15:0]   _zz_6487;
  wire       [15:0]   _zz_6488;
  wire       [15:0]   _zz_6489;
  wire       [15:0]   _zz_6490;
  wire       [15:0]   _zz_6491;
  wire       [15:0]   _zz_6492;
  wire       [15:0]   _zz_6493;
  wire       [15:0]   _zz_6494;
  wire       [15:0]   _zz_6495;
  wire       [15:0]   _zz_6496;
  wire       [31:0]   _zz_6497;
  wire       [31:0]   _zz_6498;
  wire       [15:0]   _zz_6499;
  wire       [31:0]   _zz_6500;
  wire       [31:0]   _zz_6501;
  wire       [15:0]   _zz_6502;
  wire       [15:0]   _zz_6503;
  wire       [15:0]   _zz_6504;
  wire       [15:0]   _zz_6505;
  wire       [15:0]   _zz_6506;
  wire       [15:0]   _zz_6507;
  wire       [15:0]   _zz_6508;
  wire       [15:0]   _zz_6509;
  wire       [15:0]   _zz_6510;
  wire       [15:0]   _zz_6511;
  wire       [15:0]   _zz_6512;
  wire       [15:0]   _zz_6513;
  wire       [15:0]   _zz_6514;
  wire       [15:0]   _zz_6515;
  wire       [15:0]   _zz_6516;
  wire       [15:0]   _zz_6517;
  wire       [15:0]   _zz_6518;
  wire       [31:0]   _zz_6519;
  wire       [31:0]   _zz_6520;
  wire       [15:0]   _zz_6521;
  wire       [31:0]   _zz_6522;
  wire       [31:0]   _zz_6523;
  wire       [15:0]   _zz_6524;
  wire       [15:0]   _zz_6525;
  wire       [15:0]   _zz_6526;
  wire       [15:0]   _zz_6527;
  wire       [15:0]   _zz_6528;
  wire       [15:0]   _zz_6529;
  wire       [15:0]   _zz_6530;
  wire       [15:0]   _zz_6531;
  wire       [15:0]   _zz_6532;
  wire       [15:0]   _zz_6533;
  wire       [15:0]   _zz_6534;
  wire       [15:0]   _zz_6535;
  wire       [15:0]   _zz_6536;
  wire       [15:0]   _zz_6537;
  wire       [15:0]   _zz_6538;
  wire       [15:0]   _zz_6539;
  wire       [15:0]   _zz_6540;
  wire       [31:0]   _zz_6541;
  wire       [31:0]   _zz_6542;
  wire       [15:0]   _zz_6543;
  wire       [31:0]   _zz_6544;
  wire       [31:0]   _zz_6545;
  wire       [15:0]   _zz_6546;
  wire       [15:0]   _zz_6547;
  wire       [15:0]   _zz_6548;
  wire       [15:0]   _zz_6549;
  wire       [15:0]   _zz_6550;
  wire       [15:0]   _zz_6551;
  wire       [15:0]   _zz_6552;
  wire       [15:0]   _zz_6553;
  wire       [15:0]   _zz_6554;
  wire       [15:0]   _zz_6555;
  wire       [15:0]   _zz_6556;
  wire       [15:0]   _zz_6557;
  wire       [15:0]   _zz_6558;
  wire       [15:0]   _zz_6559;
  wire       [15:0]   _zz_6560;
  wire       [15:0]   _zz_6561;
  wire       [15:0]   _zz_6562;
  wire       [31:0]   _zz_6563;
  wire       [31:0]   _zz_6564;
  wire       [15:0]   _zz_6565;
  wire       [31:0]   _zz_6566;
  wire       [31:0]   _zz_6567;
  wire       [15:0]   _zz_6568;
  wire       [15:0]   _zz_6569;
  wire       [15:0]   _zz_6570;
  wire       [15:0]   _zz_6571;
  wire       [15:0]   _zz_6572;
  wire       [15:0]   _zz_6573;
  wire       [15:0]   _zz_6574;
  wire       [15:0]   _zz_6575;
  wire       [15:0]   _zz_6576;
  wire       [15:0]   _zz_6577;
  wire       [15:0]   _zz_6578;
  wire       [15:0]   _zz_6579;
  wire       [15:0]   _zz_6580;
  wire       [15:0]   _zz_6581;
  wire       [15:0]   _zz_6582;
  wire       [15:0]   _zz_6583;
  wire       [15:0]   _zz_6584;
  wire       [31:0]   _zz_6585;
  wire       [31:0]   _zz_6586;
  wire       [15:0]   _zz_6587;
  wire       [31:0]   _zz_6588;
  wire       [31:0]   _zz_6589;
  wire       [15:0]   _zz_6590;
  wire       [15:0]   _zz_6591;
  wire       [15:0]   _zz_6592;
  wire       [15:0]   _zz_6593;
  wire       [15:0]   _zz_6594;
  wire       [15:0]   _zz_6595;
  wire       [15:0]   _zz_6596;
  wire       [15:0]   _zz_6597;
  wire       [15:0]   _zz_6598;
  wire       [15:0]   _zz_6599;
  wire       [15:0]   _zz_6600;
  wire       [15:0]   _zz_6601;
  wire       [15:0]   _zz_6602;
  wire       [15:0]   _zz_6603;
  wire       [15:0]   _zz_6604;
  wire       [15:0]   _zz_6605;
  wire       [15:0]   _zz_6606;
  wire       [31:0]   _zz_6607;
  wire       [31:0]   _zz_6608;
  wire       [15:0]   _zz_6609;
  wire       [31:0]   _zz_6610;
  wire       [31:0]   _zz_6611;
  wire       [15:0]   _zz_6612;
  wire       [15:0]   _zz_6613;
  wire       [15:0]   _zz_6614;
  wire       [15:0]   _zz_6615;
  wire       [15:0]   _zz_6616;
  wire       [15:0]   _zz_6617;
  wire       [15:0]   _zz_6618;
  wire       [15:0]   _zz_6619;
  wire       [15:0]   _zz_6620;
  wire       [15:0]   _zz_6621;
  wire       [15:0]   _zz_6622;
  wire       [15:0]   _zz_6623;
  wire       [15:0]   _zz_6624;
  wire       [15:0]   _zz_6625;
  wire       [15:0]   _zz_6626;
  wire       [15:0]   _zz_6627;
  wire       [15:0]   _zz_6628;
  wire       [31:0]   _zz_6629;
  wire       [31:0]   _zz_6630;
  wire       [15:0]   _zz_6631;
  wire       [31:0]   _zz_6632;
  wire       [31:0]   _zz_6633;
  wire       [15:0]   _zz_6634;
  wire       [15:0]   _zz_6635;
  wire       [15:0]   _zz_6636;
  wire       [15:0]   _zz_6637;
  wire       [15:0]   _zz_6638;
  wire       [15:0]   _zz_6639;
  wire       [15:0]   _zz_6640;
  wire       [15:0]   _zz_6641;
  wire       [15:0]   _zz_6642;
  wire       [15:0]   _zz_6643;
  wire       [15:0]   _zz_6644;
  wire       [15:0]   _zz_6645;
  wire       [15:0]   _zz_6646;
  wire       [15:0]   _zz_6647;
  wire       [15:0]   _zz_6648;
  wire       [15:0]   _zz_6649;
  wire       [15:0]   _zz_6650;
  wire       [31:0]   _zz_6651;
  wire       [31:0]   _zz_6652;
  wire       [15:0]   _zz_6653;
  wire       [31:0]   _zz_6654;
  wire       [31:0]   _zz_6655;
  wire       [15:0]   _zz_6656;
  wire       [15:0]   _zz_6657;
  wire       [15:0]   _zz_6658;
  wire       [15:0]   _zz_6659;
  wire       [15:0]   _zz_6660;
  wire       [15:0]   _zz_6661;
  wire       [15:0]   _zz_6662;
  wire       [15:0]   _zz_6663;
  wire       [15:0]   _zz_6664;
  wire       [15:0]   _zz_6665;
  wire       [15:0]   _zz_6666;
  wire       [15:0]   _zz_6667;
  wire       [15:0]   _zz_6668;
  wire       [15:0]   _zz_6669;
  wire       [15:0]   _zz_6670;
  wire       [15:0]   _zz_6671;
  wire       [15:0]   _zz_6672;
  wire       [31:0]   _zz_6673;
  wire       [31:0]   _zz_6674;
  wire       [15:0]   _zz_6675;
  wire       [31:0]   _zz_6676;
  wire       [31:0]   _zz_6677;
  wire       [15:0]   _zz_6678;
  wire       [15:0]   _zz_6679;
  wire       [15:0]   _zz_6680;
  wire       [15:0]   _zz_6681;
  wire       [15:0]   _zz_6682;
  wire       [15:0]   _zz_6683;
  wire       [15:0]   _zz_6684;
  wire       [15:0]   _zz_6685;
  wire       [15:0]   _zz_6686;
  wire       [15:0]   _zz_6687;
  wire       [15:0]   _zz_6688;
  wire       [15:0]   _zz_6689;
  wire       [15:0]   _zz_6690;
  wire       [15:0]   _zz_6691;
  wire       [15:0]   _zz_6692;
  wire       [15:0]   _zz_6693;
  wire       [15:0]   _zz_6694;
  wire       [31:0]   _zz_6695;
  wire       [31:0]   _zz_6696;
  wire       [15:0]   _zz_6697;
  wire       [31:0]   _zz_6698;
  wire       [31:0]   _zz_6699;
  wire       [15:0]   _zz_6700;
  wire       [15:0]   _zz_6701;
  wire       [15:0]   _zz_6702;
  wire       [15:0]   _zz_6703;
  wire       [15:0]   _zz_6704;
  wire       [15:0]   _zz_6705;
  wire       [15:0]   _zz_6706;
  wire       [15:0]   _zz_6707;
  wire       [15:0]   _zz_6708;
  wire       [15:0]   _zz_6709;
  wire       [15:0]   _zz_6710;
  wire       [15:0]   _zz_6711;
  wire       [15:0]   _zz_6712;
  wire       [15:0]   _zz_6713;
  wire       [15:0]   _zz_6714;
  wire       [15:0]   _zz_6715;
  wire       [15:0]   _zz_6716;
  wire       [31:0]   _zz_6717;
  wire       [31:0]   _zz_6718;
  wire       [15:0]   _zz_6719;
  wire       [31:0]   _zz_6720;
  wire       [31:0]   _zz_6721;
  wire       [15:0]   _zz_6722;
  wire       [15:0]   _zz_6723;
  wire       [15:0]   _zz_6724;
  wire       [15:0]   _zz_6725;
  wire       [15:0]   _zz_6726;
  wire       [15:0]   _zz_6727;
  wire       [15:0]   _zz_6728;
  wire       [15:0]   _zz_6729;
  wire       [15:0]   _zz_6730;
  wire       [15:0]   _zz_6731;
  wire       [15:0]   _zz_6732;
  wire       [15:0]   _zz_6733;
  wire       [15:0]   _zz_6734;
  wire       [15:0]   _zz_6735;
  wire       [15:0]   _zz_6736;
  wire       [15:0]   _zz_6737;
  wire       [15:0]   _zz_6738;
  wire       [31:0]   _zz_6739;
  wire       [31:0]   _zz_6740;
  wire       [15:0]   _zz_6741;
  wire       [31:0]   _zz_6742;
  wire       [31:0]   _zz_6743;
  wire       [15:0]   _zz_6744;
  wire       [15:0]   _zz_6745;
  wire       [15:0]   _zz_6746;
  wire       [15:0]   _zz_6747;
  wire       [15:0]   _zz_6748;
  wire       [15:0]   _zz_6749;
  wire       [15:0]   _zz_6750;
  wire       [15:0]   _zz_6751;
  wire       [15:0]   _zz_6752;
  wire       [15:0]   _zz_6753;
  wire       [15:0]   _zz_6754;
  wire       [15:0]   _zz_6755;
  wire       [15:0]   _zz_6756;
  wire       [15:0]   _zz_6757;
  wire       [15:0]   _zz_6758;
  wire       [15:0]   _zz_6759;
  wire       [15:0]   _zz_6760;
  wire       [31:0]   _zz_6761;
  wire       [31:0]   _zz_6762;
  wire       [15:0]   _zz_6763;
  wire       [31:0]   _zz_6764;
  wire       [31:0]   _zz_6765;
  wire       [15:0]   _zz_6766;
  wire       [15:0]   _zz_6767;
  wire       [15:0]   _zz_6768;
  wire       [15:0]   _zz_6769;
  wire       [15:0]   _zz_6770;
  wire       [15:0]   _zz_6771;
  wire       [15:0]   _zz_6772;
  wire       [15:0]   _zz_6773;
  wire       [15:0]   _zz_6774;
  wire       [15:0]   _zz_6775;
  wire       [15:0]   _zz_6776;
  wire       [15:0]   _zz_6777;
  wire       [15:0]   _zz_6778;
  wire       [15:0]   _zz_6779;
  wire       [15:0]   _zz_6780;
  wire       [15:0]   _zz_6781;
  wire       [15:0]   _zz_6782;
  wire       [31:0]   _zz_6783;
  wire       [31:0]   _zz_6784;
  wire       [15:0]   _zz_6785;
  wire       [31:0]   _zz_6786;
  wire       [31:0]   _zz_6787;
  wire       [15:0]   _zz_6788;
  wire       [15:0]   _zz_6789;
  wire       [15:0]   _zz_6790;
  wire       [15:0]   _zz_6791;
  wire       [15:0]   _zz_6792;
  wire       [15:0]   _zz_6793;
  wire       [15:0]   _zz_6794;
  wire       [15:0]   _zz_6795;
  wire       [15:0]   _zz_6796;
  wire       [15:0]   _zz_6797;
  wire       [15:0]   _zz_6798;
  wire       [15:0]   _zz_6799;
  wire       [15:0]   _zz_6800;
  wire       [15:0]   _zz_6801;
  wire       [15:0]   _zz_6802;
  wire       [15:0]   _zz_6803;
  wire       [15:0]   _zz_6804;
  wire       [31:0]   _zz_6805;
  wire       [31:0]   _zz_6806;
  wire       [15:0]   _zz_6807;
  wire       [31:0]   _zz_6808;
  wire       [31:0]   _zz_6809;
  wire       [15:0]   _zz_6810;
  wire       [15:0]   _zz_6811;
  wire       [15:0]   _zz_6812;
  wire       [15:0]   _zz_6813;
  wire       [15:0]   _zz_6814;
  wire       [15:0]   _zz_6815;
  wire       [15:0]   _zz_6816;
  wire       [15:0]   _zz_6817;
  wire       [15:0]   _zz_6818;
  wire       [15:0]   _zz_6819;
  wire       [15:0]   _zz_6820;
  wire       [15:0]   _zz_6821;
  wire       [15:0]   _zz_6822;
  wire       [15:0]   _zz_6823;
  wire       [15:0]   _zz_6824;
  wire       [15:0]   _zz_6825;
  wire       [15:0]   _zz_6826;
  wire       [31:0]   _zz_6827;
  wire       [31:0]   _zz_6828;
  wire       [15:0]   _zz_6829;
  wire       [31:0]   _zz_6830;
  wire       [31:0]   _zz_6831;
  wire       [15:0]   _zz_6832;
  wire       [15:0]   _zz_6833;
  wire       [15:0]   _zz_6834;
  wire       [15:0]   _zz_6835;
  wire       [15:0]   _zz_6836;
  wire       [15:0]   _zz_6837;
  wire       [15:0]   _zz_6838;
  wire       [15:0]   _zz_6839;
  wire       [15:0]   _zz_6840;
  wire       [15:0]   _zz_6841;
  wire       [15:0]   _zz_6842;
  wire       [15:0]   _zz_6843;
  wire       [15:0]   _zz_6844;
  wire       [15:0]   _zz_6845;
  wire       [15:0]   _zz_6846;
  wire       [15:0]   _zz_6847;
  wire       [15:0]   _zz_6848;
  wire       [31:0]   _zz_6849;
  wire       [31:0]   _zz_6850;
  wire       [15:0]   _zz_6851;
  wire       [31:0]   _zz_6852;
  wire       [31:0]   _zz_6853;
  wire       [15:0]   _zz_6854;
  wire       [15:0]   _zz_6855;
  wire       [15:0]   _zz_6856;
  wire       [15:0]   _zz_6857;
  wire       [15:0]   _zz_6858;
  wire       [15:0]   _zz_6859;
  wire       [15:0]   _zz_6860;
  wire       [15:0]   _zz_6861;
  wire       [15:0]   _zz_6862;
  wire       [15:0]   _zz_6863;
  wire       [15:0]   _zz_6864;
  wire       [15:0]   _zz_6865;
  wire       [15:0]   _zz_6866;
  wire       [15:0]   _zz_6867;
  wire       [15:0]   _zz_6868;
  wire       [15:0]   _zz_6869;
  wire       [15:0]   _zz_6870;
  wire       [31:0]   _zz_6871;
  wire       [31:0]   _zz_6872;
  wire       [15:0]   _zz_6873;
  wire       [31:0]   _zz_6874;
  wire       [31:0]   _zz_6875;
  wire       [15:0]   _zz_6876;
  wire       [15:0]   _zz_6877;
  wire       [15:0]   _zz_6878;
  wire       [15:0]   _zz_6879;
  wire       [15:0]   _zz_6880;
  wire       [15:0]   _zz_6881;
  wire       [15:0]   _zz_6882;
  wire       [15:0]   _zz_6883;
  wire       [15:0]   _zz_6884;
  wire       [15:0]   _zz_6885;
  wire       [15:0]   _zz_6886;
  wire       [15:0]   _zz_6887;
  wire       [15:0]   _zz_6888;
  wire       [15:0]   _zz_6889;
  wire       [15:0]   _zz_6890;
  wire       [15:0]   _zz_6891;
  wire       [15:0]   _zz_6892;
  wire       [31:0]   _zz_6893;
  wire       [31:0]   _zz_6894;
  wire       [15:0]   _zz_6895;
  wire       [31:0]   _zz_6896;
  wire       [31:0]   _zz_6897;
  wire       [15:0]   _zz_6898;
  wire       [15:0]   _zz_6899;
  wire       [15:0]   _zz_6900;
  wire       [15:0]   _zz_6901;
  wire       [15:0]   _zz_6902;
  wire       [15:0]   _zz_6903;
  wire       [15:0]   _zz_6904;
  wire       [15:0]   _zz_6905;
  wire       [15:0]   _zz_6906;
  wire       [15:0]   _zz_6907;
  wire       [15:0]   _zz_6908;
  wire       [15:0]   _zz_6909;
  wire       [15:0]   _zz_6910;
  wire       [15:0]   _zz_6911;
  wire       [15:0]   _zz_6912;
  wire       [15:0]   _zz_6913;
  wire       [15:0]   _zz_6914;
  wire       [31:0]   _zz_6915;
  wire       [31:0]   _zz_6916;
  wire       [15:0]   _zz_6917;
  wire       [31:0]   _zz_6918;
  wire       [31:0]   _zz_6919;
  wire       [15:0]   _zz_6920;
  wire       [15:0]   _zz_6921;
  wire       [15:0]   _zz_6922;
  wire       [15:0]   _zz_6923;
  wire       [15:0]   _zz_6924;
  wire       [15:0]   _zz_6925;
  wire       [15:0]   _zz_6926;
  wire       [15:0]   _zz_6927;
  wire       [15:0]   _zz_6928;
  wire       [15:0]   _zz_6929;
  wire       [15:0]   _zz_6930;
  wire       [15:0]   _zz_6931;
  wire       [15:0]   _zz_6932;
  wire       [15:0]   _zz_6933;
  wire       [15:0]   _zz_6934;
  wire       [15:0]   _zz_6935;
  wire       [15:0]   _zz_6936;
  wire       [31:0]   _zz_6937;
  wire       [31:0]   _zz_6938;
  wire       [15:0]   _zz_6939;
  wire       [31:0]   _zz_6940;
  wire       [31:0]   _zz_6941;
  wire       [15:0]   _zz_6942;
  wire       [15:0]   _zz_6943;
  wire       [15:0]   _zz_6944;
  wire       [15:0]   _zz_6945;
  wire       [15:0]   _zz_6946;
  wire       [15:0]   _zz_6947;
  wire       [15:0]   _zz_6948;
  wire       [15:0]   _zz_6949;
  wire       [15:0]   _zz_6950;
  wire       [15:0]   _zz_6951;
  wire       [15:0]   _zz_6952;
  wire       [15:0]   _zz_6953;
  wire       [15:0]   _zz_6954;
  wire       [15:0]   _zz_6955;
  wire       [15:0]   _zz_6956;
  wire       [15:0]   _zz_6957;
  wire       [15:0]   _zz_6958;
  wire       [31:0]   _zz_6959;
  wire       [31:0]   _zz_6960;
  wire       [15:0]   _zz_6961;
  wire       [31:0]   _zz_6962;
  wire       [31:0]   _zz_6963;
  wire       [15:0]   _zz_6964;
  wire       [15:0]   _zz_6965;
  wire       [15:0]   _zz_6966;
  wire       [15:0]   _zz_6967;
  wire       [15:0]   _zz_6968;
  wire       [15:0]   _zz_6969;
  wire       [15:0]   _zz_6970;
  wire       [15:0]   _zz_6971;
  wire       [15:0]   _zz_6972;
  wire       [15:0]   _zz_6973;
  wire       [15:0]   _zz_6974;
  wire       [15:0]   _zz_6975;
  wire       [15:0]   _zz_6976;
  wire       [15:0]   _zz_6977;
  wire       [15:0]   _zz_6978;
  wire       [15:0]   _zz_6979;
  wire       [15:0]   _zz_6980;
  wire       [31:0]   _zz_6981;
  wire       [31:0]   _zz_6982;
  wire       [15:0]   _zz_6983;
  wire       [31:0]   _zz_6984;
  wire       [31:0]   _zz_6985;
  wire       [15:0]   _zz_6986;
  wire       [15:0]   _zz_6987;
  wire       [15:0]   _zz_6988;
  wire       [15:0]   _zz_6989;
  wire       [15:0]   _zz_6990;
  wire       [15:0]   _zz_6991;
  wire       [15:0]   _zz_6992;
  wire       [15:0]   _zz_6993;
  wire       [15:0]   _zz_6994;
  wire       [15:0]   _zz_6995;
  wire       [15:0]   _zz_6996;
  wire       [15:0]   _zz_6997;
  wire       [15:0]   _zz_6998;
  wire       [15:0]   _zz_6999;
  wire       [15:0]   _zz_7000;
  wire       [15:0]   _zz_7001;
  wire       [15:0]   _zz_7002;
  wire       [31:0]   _zz_7003;
  wire       [31:0]   _zz_7004;
  wire       [15:0]   _zz_7005;
  wire       [31:0]   _zz_7006;
  wire       [31:0]   _zz_7007;
  wire       [15:0]   _zz_7008;
  wire       [15:0]   _zz_7009;
  wire       [15:0]   _zz_7010;
  wire       [15:0]   _zz_7011;
  wire       [15:0]   _zz_7012;
  wire       [15:0]   _zz_7013;
  wire       [15:0]   _zz_7014;
  wire       [15:0]   _zz_7015;
  wire       [15:0]   _zz_7016;
  wire       [15:0]   _zz_7017;
  wire       [15:0]   _zz_7018;
  wire       [15:0]   _zz_7019;
  wire       [15:0]   _zz_7020;
  wire       [15:0]   _zz_7021;
  wire       [15:0]   _zz_7022;
  wire       [15:0]   _zz_7023;
  wire       [15:0]   _zz_7024;
  wire       [31:0]   _zz_7025;
  wire       [31:0]   _zz_7026;
  wire       [15:0]   _zz_7027;
  wire       [31:0]   _zz_7028;
  wire       [31:0]   _zz_7029;
  wire       [15:0]   _zz_7030;
  wire       [15:0]   _zz_7031;
  wire       [15:0]   _zz_7032;
  wire       [15:0]   _zz_7033;
  wire       [15:0]   _zz_7034;
  wire       [15:0]   _zz_7035;
  wire       [15:0]   _zz_7036;
  wire       [15:0]   _zz_7037;
  wire       [15:0]   _zz_7038;
  wire       [15:0]   _zz_7039;
  wire       [15:0]   _zz_7040;
  wire       [15:0]   _zz_7041;
  wire       [15:0]   _zz_7042;
  wire       [15:0]   _zz_7043;
  wire       [15:0]   _zz_7044;
  wire       [15:0]   _zz_7045;
  wire       [15:0]   _zz_7046;
  wire       [31:0]   _zz_7047;
  wire       [31:0]   _zz_7048;
  wire       [15:0]   _zz_7049;
  wire       [31:0]   _zz_7050;
  wire       [31:0]   _zz_7051;
  wire       [15:0]   _zz_7052;
  wire       [15:0]   _zz_7053;
  wire       [15:0]   _zz_7054;
  wire       [15:0]   _zz_7055;
  wire       [15:0]   _zz_7056;
  wire       [15:0]   _zz_7057;
  wire       [15:0]   _zz_7058;
  wire       [15:0]   _zz_7059;
  wire       [15:0]   _zz_7060;
  wire       [15:0]   _zz_7061;
  wire       [15:0]   _zz_7062;
  wire       [15:0]   _zz_7063;
  wire       [15:0]   _zz_7064;
  wire       [15:0]   _zz_7065;
  wire       [15:0]   _zz_7066;
  wire       [15:0]   _zz_7067;
  wire       [15:0]   _zz_7068;
  wire       [31:0]   _zz_7069;
  wire       [31:0]   _zz_7070;
  wire       [15:0]   _zz_7071;
  wire       [31:0]   _zz_7072;
  wire       [31:0]   _zz_7073;
  wire       [15:0]   _zz_7074;
  wire       [15:0]   _zz_7075;
  wire       [15:0]   _zz_7076;
  wire       [15:0]   _zz_7077;
  wire       [15:0]   _zz_7078;
  wire       [15:0]   _zz_7079;
  wire       [15:0]   _zz_7080;
  wire       [15:0]   _zz_7081;
  wire       [15:0]   _zz_7082;
  wire       [15:0]   _zz_7083;
  wire       [15:0]   _zz_7084;
  wire       [15:0]   _zz_7085;
  wire       [15:0]   _zz_7086;
  wire       [15:0]   _zz_7087;
  wire       [15:0]   _zz_7088;
  wire       [15:0]   _zz_7089;
  wire       [15:0]   _zz_7090;
  wire       [31:0]   _zz_7091;
  wire       [31:0]   _zz_7092;
  wire       [15:0]   _zz_7093;
  wire       [31:0]   _zz_7094;
  wire       [31:0]   _zz_7095;
  wire       [15:0]   _zz_7096;
  wire       [15:0]   _zz_7097;
  wire       [15:0]   _zz_7098;
  wire       [15:0]   _zz_7099;
  wire       [15:0]   _zz_7100;
  wire       [15:0]   _zz_7101;
  wire       [15:0]   _zz_7102;
  wire       [15:0]   _zz_7103;
  wire       [15:0]   _zz_7104;
  wire       [15:0]   _zz_7105;
  wire       [15:0]   _zz_7106;
  wire       [15:0]   _zz_7107;
  wire       [15:0]   _zz_7108;
  wire       [15:0]   _zz_7109;
  wire       [15:0]   _zz_7110;
  wire       [15:0]   _zz_7111;
  wire       [15:0]   _zz_7112;
  wire       [31:0]   _zz_7113;
  wire       [31:0]   _zz_7114;
  wire       [15:0]   _zz_7115;
  wire       [31:0]   _zz_7116;
  wire       [31:0]   _zz_7117;
  wire       [15:0]   _zz_7118;
  wire       [15:0]   _zz_7119;
  wire       [15:0]   _zz_7120;
  wire       [15:0]   _zz_7121;
  wire       [15:0]   _zz_7122;
  wire       [15:0]   _zz_7123;
  wire       [15:0]   _zz_7124;
  wire       [15:0]   _zz_7125;
  wire       [15:0]   _zz_7126;
  wire       [15:0]   _zz_7127;
  wire       [15:0]   _zz_7128;
  wire       [15:0]   _zz_7129;
  wire       [15:0]   _zz_7130;
  wire       [15:0]   _zz_7131;
  wire       [15:0]   _zz_7132;
  wire       [15:0]   _zz_7133;
  wire       [15:0]   _zz_7134;
  wire       [31:0]   _zz_7135;
  wire       [31:0]   _zz_7136;
  wire       [15:0]   _zz_7137;
  wire       [31:0]   _zz_7138;
  wire       [31:0]   _zz_7139;
  wire       [15:0]   _zz_7140;
  wire       [15:0]   _zz_7141;
  wire       [15:0]   _zz_7142;
  wire       [15:0]   _zz_7143;
  wire       [15:0]   _zz_7144;
  wire       [15:0]   _zz_7145;
  wire       [15:0]   _zz_7146;
  wire       [15:0]   _zz_7147;
  wire       [15:0]   _zz_7148;
  wire       [15:0]   _zz_7149;
  wire       [15:0]   _zz_7150;
  wire       [15:0]   _zz_7151;
  wire       [15:0]   _zz_7152;
  wire       [15:0]   _zz_7153;
  wire       [15:0]   _zz_7154;
  wire       [15:0]   _zz_7155;
  wire       [15:0]   _zz_7156;
  wire       [31:0]   _zz_7157;
  wire       [31:0]   _zz_7158;
  wire       [15:0]   _zz_7159;
  wire       [31:0]   _zz_7160;
  wire       [31:0]   _zz_7161;
  wire       [15:0]   _zz_7162;
  wire       [15:0]   _zz_7163;
  wire       [15:0]   _zz_7164;
  wire       [15:0]   _zz_7165;
  wire       [15:0]   _zz_7166;
  wire       [15:0]   _zz_7167;
  wire       [15:0]   _zz_7168;
  wire       [15:0]   _zz_7169;
  wire       [15:0]   _zz_7170;
  wire       [15:0]   _zz_7171;
  wire       [15:0]   _zz_7172;
  wire       [15:0]   _zz_7173;
  wire       [15:0]   _zz_7174;
  wire       [15:0]   _zz_7175;
  wire       [15:0]   _zz_7176;
  wire       [15:0]   _zz_7177;
  wire       [15:0]   _zz_7178;
  wire       [31:0]   _zz_7179;
  wire       [31:0]   _zz_7180;
  wire       [15:0]   _zz_7181;
  wire       [31:0]   _zz_7182;
  wire       [31:0]   _zz_7183;
  wire       [15:0]   _zz_7184;
  wire       [15:0]   _zz_7185;
  wire       [15:0]   _zz_7186;
  wire       [15:0]   _zz_7187;
  wire       [15:0]   _zz_7188;
  wire       [15:0]   _zz_7189;
  wire       [15:0]   _zz_7190;
  wire       [15:0]   _zz_7191;
  wire       [15:0]   _zz_7192;
  wire       [15:0]   _zz_7193;
  wire       [15:0]   _zz_7194;
  wire       [15:0]   _zz_7195;
  wire       [15:0]   _zz_7196;
  wire       [15:0]   _zz_7197;
  wire       [15:0]   _zz_7198;
  wire       [15:0]   _zz_7199;
  wire       [15:0]   _zz_7200;
  wire       [31:0]   _zz_7201;
  wire       [31:0]   _zz_7202;
  wire       [15:0]   _zz_7203;
  wire       [31:0]   _zz_7204;
  wire       [31:0]   _zz_7205;
  wire       [15:0]   _zz_7206;
  wire       [15:0]   _zz_7207;
  wire       [15:0]   _zz_7208;
  wire       [15:0]   _zz_7209;
  wire       [15:0]   _zz_7210;
  wire       [15:0]   _zz_7211;
  wire       [15:0]   _zz_7212;
  wire       [15:0]   _zz_7213;
  wire       [15:0]   _zz_7214;
  wire       [15:0]   _zz_7215;
  wire       [15:0]   _zz_7216;
  wire       [15:0]   _zz_7217;
  wire       [15:0]   _zz_7218;
  wire       [15:0]   _zz_7219;
  wire       [15:0]   _zz_7220;
  wire       [15:0]   _zz_7221;
  wire       [15:0]   _zz_7222;
  wire       [31:0]   _zz_7223;
  wire       [31:0]   _zz_7224;
  wire       [15:0]   _zz_7225;
  wire       [31:0]   _zz_7226;
  wire       [31:0]   _zz_7227;
  wire       [15:0]   _zz_7228;
  wire       [15:0]   _zz_7229;
  wire       [15:0]   _zz_7230;
  wire       [15:0]   _zz_7231;
  wire       [15:0]   _zz_7232;
  wire       [15:0]   _zz_7233;
  wire       [15:0]   _zz_7234;
  wire       [15:0]   _zz_7235;
  wire       [15:0]   _zz_7236;
  wire       [15:0]   _zz_7237;
  wire       [15:0]   _zz_7238;
  wire       [15:0]   _zz_7239;
  wire       [15:0]   _zz_7240;
  wire       [15:0]   _zz_7241;
  wire       [15:0]   _zz_7242;
  wire       [15:0]   _zz_7243;
  wire       [15:0]   _zz_7244;
  wire       [31:0]   _zz_7245;
  wire       [31:0]   _zz_7246;
  wire       [15:0]   _zz_7247;
  wire       [31:0]   _zz_7248;
  wire       [31:0]   _zz_7249;
  wire       [15:0]   _zz_7250;
  wire       [15:0]   _zz_7251;
  wire       [15:0]   _zz_7252;
  wire       [15:0]   _zz_7253;
  wire       [15:0]   _zz_7254;
  wire       [15:0]   _zz_7255;
  wire       [15:0]   _zz_7256;
  wire       [15:0]   _zz_7257;
  wire       [15:0]   _zz_7258;
  wire       [15:0]   _zz_7259;
  wire       [15:0]   _zz_7260;
  wire       [15:0]   _zz_7261;
  wire       [15:0]   _zz_7262;
  wire       [15:0]   _zz_7263;
  wire       [15:0]   _zz_7264;
  wire       [15:0]   _zz_7265;
  wire       [15:0]   _zz_7266;
  wire       [31:0]   _zz_7267;
  wire       [31:0]   _zz_7268;
  wire       [15:0]   _zz_7269;
  wire       [31:0]   _zz_7270;
  wire       [31:0]   _zz_7271;
  wire       [15:0]   _zz_7272;
  wire       [15:0]   _zz_7273;
  wire       [15:0]   _zz_7274;
  wire       [15:0]   _zz_7275;
  wire       [15:0]   _zz_7276;
  wire       [15:0]   _zz_7277;
  wire       [15:0]   _zz_7278;
  wire       [15:0]   _zz_7279;
  wire       [15:0]   _zz_7280;
  wire       [15:0]   _zz_7281;
  wire       [15:0]   _zz_7282;
  wire       [15:0]   _zz_7283;
  wire       [15:0]   _zz_7284;
  wire       [15:0]   _zz_7285;
  wire       [15:0]   _zz_7286;
  wire       [15:0]   _zz_7287;
  wire       [15:0]   _zz_7288;
  wire       [31:0]   _zz_7289;
  wire       [31:0]   _zz_7290;
  wire       [15:0]   _zz_7291;
  wire       [31:0]   _zz_7292;
  wire       [31:0]   _zz_7293;
  wire       [15:0]   _zz_7294;
  wire       [15:0]   _zz_7295;
  wire       [15:0]   _zz_7296;
  wire       [15:0]   _zz_7297;
  wire       [15:0]   _zz_7298;
  wire       [15:0]   _zz_7299;
  wire       [15:0]   _zz_7300;
  wire       [15:0]   _zz_7301;
  wire       [15:0]   _zz_7302;
  wire       [15:0]   _zz_7303;
  wire       [15:0]   _zz_7304;
  wire       [15:0]   _zz_7305;
  wire       [15:0]   _zz_7306;
  wire       [15:0]   _zz_7307;
  wire       [15:0]   _zz_7308;
  wire       [15:0]   _zz_7309;
  wire       [15:0]   _zz_7310;
  wire       [31:0]   _zz_7311;
  wire       [31:0]   _zz_7312;
  wire       [15:0]   _zz_7313;
  wire       [31:0]   _zz_7314;
  wire       [31:0]   _zz_7315;
  wire       [15:0]   _zz_7316;
  wire       [15:0]   _zz_7317;
  wire       [15:0]   _zz_7318;
  wire       [15:0]   _zz_7319;
  wire       [15:0]   _zz_7320;
  wire       [15:0]   _zz_7321;
  wire       [15:0]   _zz_7322;
  wire       [15:0]   _zz_7323;
  wire       [15:0]   _zz_7324;
  wire       [15:0]   _zz_7325;
  wire       [15:0]   _zz_7326;
  wire       [15:0]   _zz_7327;
  wire       [15:0]   _zz_7328;
  wire       [15:0]   _zz_7329;
  wire       [15:0]   _zz_7330;
  wire       [15:0]   _zz_7331;
  wire       [15:0]   _zz_7332;
  wire       [31:0]   _zz_7333;
  wire       [31:0]   _zz_7334;
  wire       [15:0]   _zz_7335;
  wire       [31:0]   _zz_7336;
  wire       [31:0]   _zz_7337;
  wire       [15:0]   _zz_7338;
  wire       [15:0]   _zz_7339;
  wire       [15:0]   _zz_7340;
  wire       [15:0]   _zz_7341;
  wire       [15:0]   _zz_7342;
  wire       [15:0]   _zz_7343;
  wire       [15:0]   _zz_7344;
  wire       [15:0]   _zz_7345;
  wire       [15:0]   _zz_7346;
  wire       [15:0]   _zz_7347;
  wire       [15:0]   _zz_7348;
  wire       [15:0]   _zz_7349;
  wire       [15:0]   _zz_7350;
  wire       [15:0]   _zz_7351;
  wire       [15:0]   _zz_7352;
  wire       [15:0]   _zz_7353;
  wire       [15:0]   _zz_7354;
  wire       [31:0]   _zz_7355;
  wire       [31:0]   _zz_7356;
  wire       [15:0]   _zz_7357;
  wire       [31:0]   _zz_7358;
  wire       [31:0]   _zz_7359;
  wire       [15:0]   _zz_7360;
  wire       [15:0]   _zz_7361;
  wire       [15:0]   _zz_7362;
  wire       [15:0]   _zz_7363;
  wire       [15:0]   _zz_7364;
  wire       [15:0]   _zz_7365;
  wire       [15:0]   _zz_7366;
  wire       [15:0]   _zz_7367;
  wire       [15:0]   _zz_7368;
  wire       [15:0]   _zz_7369;
  wire       [15:0]   _zz_7370;
  wire       [15:0]   _zz_7371;
  wire       [15:0]   _zz_7372;
  wire       [15:0]   _zz_7373;
  wire       [15:0]   _zz_7374;
  wire       [15:0]   _zz_7375;
  wire       [15:0]   _zz_7376;
  wire       [31:0]   _zz_7377;
  wire       [31:0]   _zz_7378;
  wire       [15:0]   _zz_7379;
  wire       [31:0]   _zz_7380;
  wire       [31:0]   _zz_7381;
  wire       [15:0]   _zz_7382;
  wire       [15:0]   _zz_7383;
  wire       [15:0]   _zz_7384;
  wire       [15:0]   _zz_7385;
  wire       [15:0]   _zz_7386;
  wire       [15:0]   _zz_7387;
  wire       [15:0]   _zz_7388;
  wire       [15:0]   _zz_7389;
  wire       [15:0]   _zz_7390;
  wire       [15:0]   _zz_7391;
  wire       [15:0]   _zz_7392;
  wire       [15:0]   _zz_7393;
  wire       [15:0]   _zz_7394;
  wire       [15:0]   _zz_7395;
  wire       [15:0]   _zz_7396;
  wire       [15:0]   _zz_7397;
  wire       [15:0]   _zz_7398;
  wire       [31:0]   _zz_7399;
  wire       [31:0]   _zz_7400;
  wire       [15:0]   _zz_7401;
  wire       [31:0]   _zz_7402;
  wire       [31:0]   _zz_7403;
  wire       [15:0]   _zz_7404;
  wire       [15:0]   _zz_7405;
  wire       [15:0]   _zz_7406;
  wire       [15:0]   _zz_7407;
  wire       [15:0]   _zz_7408;
  wire       [15:0]   _zz_7409;
  wire       [15:0]   _zz_7410;
  wire       [15:0]   _zz_7411;
  wire       [15:0]   _zz_7412;
  wire       [15:0]   _zz_7413;
  wire       [15:0]   _zz_7414;
  wire       [15:0]   _zz_7415;
  wire       [15:0]   _zz_7416;
  wire       [15:0]   _zz_7417;
  wire       [15:0]   _zz_7418;
  wire       [15:0]   _zz_7419;
  wire       [15:0]   _zz_7420;
  wire       [31:0]   _zz_7421;
  wire       [31:0]   _zz_7422;
  wire       [15:0]   _zz_7423;
  wire       [31:0]   _zz_7424;
  wire       [31:0]   _zz_7425;
  wire       [15:0]   _zz_7426;
  wire       [15:0]   _zz_7427;
  wire       [15:0]   _zz_7428;
  wire       [15:0]   _zz_7429;
  wire       [15:0]   _zz_7430;
  wire       [15:0]   _zz_7431;
  wire       [15:0]   _zz_7432;
  wire       [15:0]   _zz_7433;
  wire       [15:0]   _zz_7434;
  wire       [15:0]   _zz_7435;
  wire       [15:0]   _zz_7436;
  wire       [15:0]   _zz_7437;
  wire       [15:0]   _zz_7438;
  wire       [15:0]   _zz_7439;
  wire       [15:0]   _zz_7440;
  wire       [15:0]   _zz_7441;
  wire       [15:0]   _zz_7442;
  wire       [31:0]   _zz_7443;
  wire       [31:0]   _zz_7444;
  wire       [15:0]   _zz_7445;
  wire       [31:0]   _zz_7446;
  wire       [31:0]   _zz_7447;
  wire       [15:0]   _zz_7448;
  wire       [15:0]   _zz_7449;
  wire       [15:0]   _zz_7450;
  wire       [15:0]   _zz_7451;
  wire       [15:0]   _zz_7452;
  wire       [15:0]   _zz_7453;
  wire       [15:0]   _zz_7454;
  wire       [15:0]   _zz_7455;
  wire       [15:0]   _zz_7456;
  wire       [15:0]   _zz_7457;
  wire       [15:0]   _zz_7458;
  wire       [15:0]   _zz_7459;
  wire       [15:0]   _zz_7460;
  wire       [15:0]   _zz_7461;
  wire       [15:0]   _zz_7462;
  wire       [15:0]   _zz_7463;
  wire       [15:0]   _zz_7464;
  wire       [31:0]   _zz_7465;
  wire       [31:0]   _zz_7466;
  wire       [15:0]   _zz_7467;
  wire       [31:0]   _zz_7468;
  wire       [31:0]   _zz_7469;
  wire       [15:0]   _zz_7470;
  wire       [15:0]   _zz_7471;
  wire       [15:0]   _zz_7472;
  wire       [15:0]   _zz_7473;
  wire       [15:0]   _zz_7474;
  wire       [15:0]   _zz_7475;
  wire       [15:0]   _zz_7476;
  wire       [15:0]   _zz_7477;
  wire       [15:0]   _zz_7478;
  wire       [15:0]   _zz_7479;
  wire       [15:0]   _zz_7480;
  wire       [15:0]   _zz_7481;
  wire       [15:0]   _zz_7482;
  wire       [15:0]   _zz_7483;
  wire       [15:0]   _zz_7484;
  wire       [15:0]   _zz_7485;
  wire       [15:0]   _zz_7486;
  wire       [31:0]   _zz_7487;
  wire       [31:0]   _zz_7488;
  wire       [15:0]   _zz_7489;
  wire       [31:0]   _zz_7490;
  wire       [31:0]   _zz_7491;
  wire       [15:0]   _zz_7492;
  wire       [15:0]   _zz_7493;
  wire       [15:0]   _zz_7494;
  wire       [15:0]   _zz_7495;
  wire       [15:0]   _zz_7496;
  wire       [15:0]   _zz_7497;
  wire       [15:0]   _zz_7498;
  wire       [15:0]   _zz_7499;
  wire       [15:0]   _zz_7500;
  wire       [15:0]   _zz_7501;
  wire       [15:0]   _zz_7502;
  wire       [15:0]   _zz_7503;
  wire       [15:0]   _zz_7504;
  wire       [15:0]   _zz_7505;
  wire       [15:0]   _zz_7506;
  wire       [15:0]   _zz_7507;
  wire       [15:0]   _zz_7508;
  wire       [31:0]   _zz_7509;
  wire       [31:0]   _zz_7510;
  wire       [15:0]   _zz_7511;
  wire       [31:0]   _zz_7512;
  wire       [31:0]   _zz_7513;
  wire       [15:0]   _zz_7514;
  wire       [15:0]   _zz_7515;
  wire       [15:0]   _zz_7516;
  wire       [15:0]   _zz_7517;
  wire       [15:0]   _zz_7518;
  wire       [15:0]   _zz_7519;
  wire       [15:0]   _zz_7520;
  wire       [15:0]   _zz_7521;
  wire       [15:0]   _zz_7522;
  wire       [15:0]   _zz_7523;
  wire       [15:0]   _zz_7524;
  wire       [15:0]   _zz_7525;
  wire       [15:0]   _zz_7526;
  wire       [15:0]   _zz_7527;
  wire       [15:0]   _zz_7528;
  wire       [15:0]   _zz_7529;
  wire       [15:0]   _zz_7530;
  wire       [31:0]   _zz_7531;
  wire       [31:0]   _zz_7532;
  wire       [15:0]   _zz_7533;
  wire       [31:0]   _zz_7534;
  wire       [31:0]   _zz_7535;
  wire       [15:0]   _zz_7536;
  wire       [15:0]   _zz_7537;
  wire       [15:0]   _zz_7538;
  wire       [15:0]   _zz_7539;
  wire       [15:0]   _zz_7540;
  wire       [15:0]   _zz_7541;
  wire       [15:0]   _zz_7542;
  wire       [15:0]   _zz_7543;
  wire       [15:0]   _zz_7544;
  wire       [15:0]   _zz_7545;
  wire       [15:0]   _zz_7546;
  wire       [15:0]   _zz_7547;
  wire       [15:0]   _zz_7548;
  wire       [15:0]   _zz_7549;
  wire       [15:0]   _zz_7550;
  wire       [15:0]   _zz_7551;
  wire       [15:0]   _zz_7552;
  wire       [31:0]   _zz_7553;
  wire       [31:0]   _zz_7554;
  wire       [15:0]   _zz_7555;
  wire       [31:0]   _zz_7556;
  wire       [31:0]   _zz_7557;
  wire       [15:0]   _zz_7558;
  wire       [15:0]   _zz_7559;
  wire       [15:0]   _zz_7560;
  wire       [15:0]   _zz_7561;
  wire       [15:0]   _zz_7562;
  wire       [15:0]   _zz_7563;
  wire       [15:0]   _zz_7564;
  wire       [15:0]   _zz_7565;
  wire       [15:0]   _zz_7566;
  wire       [15:0]   _zz_7567;
  wire       [15:0]   _zz_7568;
  wire       [15:0]   _zz_7569;
  wire       [15:0]   _zz_7570;
  wire       [15:0]   _zz_7571;
  wire       [15:0]   _zz_7572;
  wire       [15:0]   _zz_7573;
  wire       [15:0]   _zz_7574;
  wire       [31:0]   _zz_7575;
  wire       [31:0]   _zz_7576;
  wire       [15:0]   _zz_7577;
  wire       [31:0]   _zz_7578;
  wire       [31:0]   _zz_7579;
  wire       [15:0]   _zz_7580;
  wire       [15:0]   _zz_7581;
  wire       [15:0]   _zz_7582;
  wire       [15:0]   _zz_7583;
  wire       [15:0]   _zz_7584;
  wire       [15:0]   _zz_7585;
  wire       [15:0]   _zz_7586;
  wire       [15:0]   _zz_7587;
  wire       [15:0]   _zz_7588;
  wire       [15:0]   _zz_7589;
  wire       [15:0]   _zz_7590;
  wire       [15:0]   _zz_7591;
  wire       [15:0]   _zz_7592;
  wire       [15:0]   _zz_7593;
  wire       [15:0]   _zz_7594;
  wire       [15:0]   _zz_7595;
  wire       [15:0]   _zz_7596;
  wire       [31:0]   _zz_7597;
  wire       [31:0]   _zz_7598;
  wire       [15:0]   _zz_7599;
  wire       [31:0]   _zz_7600;
  wire       [31:0]   _zz_7601;
  wire       [15:0]   _zz_7602;
  wire       [15:0]   _zz_7603;
  wire       [15:0]   _zz_7604;
  wire       [15:0]   _zz_7605;
  wire       [15:0]   _zz_7606;
  wire       [15:0]   _zz_7607;
  wire       [15:0]   _zz_7608;
  wire       [15:0]   _zz_7609;
  wire       [15:0]   _zz_7610;
  wire       [15:0]   _zz_7611;
  wire       [15:0]   _zz_7612;
  wire       [15:0]   _zz_7613;
  wire       [15:0]   _zz_7614;
  wire       [15:0]   _zz_7615;
  wire       [15:0]   _zz_7616;
  wire       [15:0]   _zz_7617;
  wire       [15:0]   _zz_7618;
  wire       [31:0]   _zz_7619;
  wire       [31:0]   _zz_7620;
  wire       [15:0]   _zz_7621;
  wire       [31:0]   _zz_7622;
  wire       [31:0]   _zz_7623;
  wire       [15:0]   _zz_7624;
  wire       [15:0]   _zz_7625;
  wire       [15:0]   _zz_7626;
  wire       [15:0]   _zz_7627;
  wire       [15:0]   _zz_7628;
  wire       [15:0]   _zz_7629;
  wire       [15:0]   _zz_7630;
  wire       [15:0]   _zz_7631;
  wire       [15:0]   _zz_7632;
  wire       [15:0]   _zz_7633;
  wire       [15:0]   _zz_7634;
  wire       [15:0]   _zz_7635;
  wire       [15:0]   _zz_7636;
  wire       [15:0]   _zz_7637;
  wire       [15:0]   _zz_7638;
  wire       [15:0]   _zz_7639;
  wire       [15:0]   _zz_7640;
  wire       [31:0]   _zz_7641;
  wire       [31:0]   _zz_7642;
  wire       [15:0]   _zz_7643;
  wire       [31:0]   _zz_7644;
  wire       [31:0]   _zz_7645;
  wire       [15:0]   _zz_7646;
  wire       [15:0]   _zz_7647;
  wire       [15:0]   _zz_7648;
  wire       [15:0]   _zz_7649;
  wire       [15:0]   _zz_7650;
  wire       [15:0]   _zz_7651;
  wire       [15:0]   _zz_7652;
  wire       [15:0]   _zz_7653;
  wire       [15:0]   _zz_7654;
  wire       [15:0]   _zz_7655;
  wire       [15:0]   _zz_7656;
  wire       [15:0]   _zz_7657;
  wire       [15:0]   _zz_7658;
  wire       [15:0]   _zz_7659;
  wire       [15:0]   _zz_7660;
  wire       [15:0]   _zz_7661;
  wire       [15:0]   _zz_7662;
  wire       [31:0]   _zz_7663;
  wire       [31:0]   _zz_7664;
  wire       [15:0]   _zz_7665;
  wire       [31:0]   _zz_7666;
  wire       [31:0]   _zz_7667;
  wire       [15:0]   _zz_7668;
  wire       [15:0]   _zz_7669;
  wire       [15:0]   _zz_7670;
  wire       [15:0]   _zz_7671;
  wire       [15:0]   _zz_7672;
  wire       [15:0]   _zz_7673;
  wire       [15:0]   _zz_7674;
  wire       [15:0]   _zz_7675;
  wire       [15:0]   _zz_7676;
  wire       [15:0]   _zz_7677;
  wire       [15:0]   _zz_7678;
  wire       [15:0]   _zz_7679;
  wire       [15:0]   _zz_7680;
  wire       [15:0]   _zz_7681;
  wire       [15:0]   _zz_7682;
  wire       [15:0]   _zz_7683;
  wire       [15:0]   _zz_7684;
  wire       [31:0]   _zz_7685;
  wire       [31:0]   _zz_7686;
  wire       [15:0]   _zz_7687;
  wire       [31:0]   _zz_7688;
  wire       [31:0]   _zz_7689;
  wire       [15:0]   _zz_7690;
  wire       [15:0]   _zz_7691;
  wire       [15:0]   _zz_7692;
  wire       [15:0]   _zz_7693;
  wire       [15:0]   _zz_7694;
  wire       [15:0]   _zz_7695;
  wire       [15:0]   _zz_7696;
  wire       [15:0]   _zz_7697;
  wire       [15:0]   _zz_7698;
  wire       [15:0]   _zz_7699;
  wire       [15:0]   _zz_7700;
  wire       [15:0]   _zz_7701;
  wire       [15:0]   _zz_7702;
  wire       [15:0]   _zz_7703;
  wire       [15:0]   _zz_7704;
  wire       [15:0]   _zz_7705;
  wire       [15:0]   _zz_7706;
  wire       [31:0]   _zz_7707;
  wire       [31:0]   _zz_7708;
  wire       [15:0]   _zz_7709;
  wire       [31:0]   _zz_7710;
  wire       [31:0]   _zz_7711;
  wire       [15:0]   _zz_7712;
  wire       [15:0]   _zz_7713;
  wire       [15:0]   _zz_7714;
  wire       [15:0]   _zz_7715;
  wire       [15:0]   _zz_7716;
  wire       [15:0]   _zz_7717;
  wire       [15:0]   _zz_7718;
  wire       [15:0]   _zz_7719;
  wire       [15:0]   _zz_7720;
  wire       [15:0]   _zz_7721;
  wire       [15:0]   _zz_7722;
  wire       [15:0]   _zz_7723;
  wire       [15:0]   _zz_7724;
  wire       [15:0]   _zz_7725;
  wire       [15:0]   _zz_7726;
  wire       [15:0]   _zz_7727;
  wire       [15:0]   _zz_7728;
  wire       [31:0]   _zz_7729;
  wire       [31:0]   _zz_7730;
  wire       [15:0]   _zz_7731;
  wire       [31:0]   _zz_7732;
  wire       [31:0]   _zz_7733;
  wire       [15:0]   _zz_7734;
  wire       [15:0]   _zz_7735;
  wire       [15:0]   _zz_7736;
  wire       [15:0]   _zz_7737;
  wire       [15:0]   _zz_7738;
  wire       [15:0]   _zz_7739;
  wire       [15:0]   _zz_7740;
  wire       [15:0]   _zz_7741;
  wire       [15:0]   _zz_7742;
  wire       [15:0]   _zz_7743;
  wire       [15:0]   _zz_7744;
  wire       [15:0]   _zz_7745;
  wire       [15:0]   _zz_7746;
  wire       [15:0]   _zz_7747;
  wire       [15:0]   _zz_7748;
  wire       [15:0]   _zz_7749;
  wire       [15:0]   _zz_7750;
  wire       [31:0]   _zz_7751;
  wire       [31:0]   _zz_7752;
  wire       [15:0]   _zz_7753;
  wire       [31:0]   _zz_7754;
  wire       [31:0]   _zz_7755;
  wire       [15:0]   _zz_7756;
  wire       [15:0]   _zz_7757;
  wire       [15:0]   _zz_7758;
  wire       [15:0]   _zz_7759;
  wire       [15:0]   _zz_7760;
  wire       [15:0]   _zz_7761;
  wire       [15:0]   _zz_7762;
  wire       [15:0]   _zz_7763;
  wire       [15:0]   _zz_7764;
  wire       [15:0]   _zz_7765;
  wire       [15:0]   _zz_7766;
  wire       [15:0]   _zz_7767;
  wire       [15:0]   _zz_7768;
  wire       [15:0]   _zz_7769;
  wire       [15:0]   _zz_7770;
  wire       [15:0]   _zz_7771;
  wire       [15:0]   _zz_7772;
  wire       [31:0]   _zz_7773;
  wire       [31:0]   _zz_7774;
  wire       [15:0]   _zz_7775;
  wire       [31:0]   _zz_7776;
  wire       [31:0]   _zz_7777;
  wire       [15:0]   _zz_7778;
  wire       [15:0]   _zz_7779;
  wire       [15:0]   _zz_7780;
  wire       [15:0]   _zz_7781;
  wire       [15:0]   _zz_7782;
  wire       [15:0]   _zz_7783;
  wire       [15:0]   _zz_7784;
  wire       [15:0]   _zz_7785;
  wire       [15:0]   _zz_7786;
  wire       [15:0]   _zz_7787;
  wire       [15:0]   _zz_7788;
  wire       [15:0]   _zz_7789;
  wire       [15:0]   _zz_7790;
  wire       [15:0]   _zz_7791;
  wire       [15:0]   _zz_7792;
  wire       [15:0]   _zz_7793;
  wire       [15:0]   _zz_7794;
  wire       [31:0]   _zz_7795;
  wire       [31:0]   _zz_7796;
  wire       [15:0]   _zz_7797;
  wire       [31:0]   _zz_7798;
  wire       [31:0]   _zz_7799;
  wire       [15:0]   _zz_7800;
  wire       [15:0]   _zz_7801;
  wire       [15:0]   _zz_7802;
  wire       [15:0]   _zz_7803;
  wire       [15:0]   _zz_7804;
  wire       [15:0]   _zz_7805;
  wire       [15:0]   _zz_7806;
  wire       [15:0]   _zz_7807;
  wire       [15:0]   _zz_7808;
  wire       [15:0]   _zz_7809;
  wire       [15:0]   _zz_7810;
  wire       [15:0]   _zz_7811;
  wire       [15:0]   _zz_7812;
  wire       [15:0]   _zz_7813;
  wire       [15:0]   _zz_7814;
  wire       [15:0]   _zz_7815;
  wire       [15:0]   _zz_7816;
  wire       [31:0]   _zz_7817;
  wire       [31:0]   _zz_7818;
  wire       [15:0]   _zz_7819;
  wire       [31:0]   _zz_7820;
  wire       [31:0]   _zz_7821;
  wire       [15:0]   _zz_7822;
  wire       [15:0]   _zz_7823;
  wire       [15:0]   _zz_7824;
  wire       [15:0]   _zz_7825;
  wire       [15:0]   _zz_7826;
  wire       [15:0]   _zz_7827;
  wire       [15:0]   _zz_7828;
  wire       [15:0]   _zz_7829;
  wire       [15:0]   _zz_7830;
  wire       [15:0]   _zz_7831;
  wire       [15:0]   _zz_7832;
  wire       [15:0]   _zz_7833;
  wire       [15:0]   _zz_7834;
  wire       [15:0]   _zz_7835;
  wire       [15:0]   _zz_7836;
  wire       [15:0]   _zz_7837;
  wire       [15:0]   _zz_7838;
  wire       [31:0]   _zz_7839;
  wire       [31:0]   _zz_7840;
  wire       [15:0]   _zz_7841;
  wire       [31:0]   _zz_7842;
  wire       [31:0]   _zz_7843;
  wire       [15:0]   _zz_7844;
  wire       [15:0]   _zz_7845;
  wire       [15:0]   _zz_7846;
  wire       [15:0]   _zz_7847;
  wire       [15:0]   _zz_7848;
  wire       [15:0]   _zz_7849;
  wire       [15:0]   _zz_7850;
  wire       [15:0]   _zz_7851;
  wire       [15:0]   _zz_7852;
  wire       [15:0]   _zz_7853;
  wire       [15:0]   _zz_7854;
  wire       [15:0]   _zz_7855;
  wire       [15:0]   _zz_7856;
  wire       [15:0]   _zz_7857;
  wire       [15:0]   _zz_7858;
  wire       [15:0]   _zz_7859;
  wire       [15:0]   _zz_7860;
  wire       [31:0]   _zz_7861;
  wire       [31:0]   _zz_7862;
  wire       [15:0]   _zz_7863;
  wire       [31:0]   _zz_7864;
  wire       [31:0]   _zz_7865;
  wire       [15:0]   _zz_7866;
  wire       [15:0]   _zz_7867;
  wire       [15:0]   _zz_7868;
  wire       [15:0]   _zz_7869;
  wire       [15:0]   _zz_7870;
  wire       [15:0]   _zz_7871;
  wire       [15:0]   _zz_7872;
  wire       [15:0]   _zz_7873;
  wire       [15:0]   _zz_7874;
  wire       [15:0]   _zz_7875;
  wire       [15:0]   _zz_7876;
  wire       [15:0]   _zz_7877;
  wire       [15:0]   _zz_7878;
  wire       [15:0]   _zz_7879;
  wire       [15:0]   _zz_7880;
  wire       [15:0]   _zz_7881;
  wire       [15:0]   _zz_7882;
  wire       [31:0]   _zz_7883;
  wire       [31:0]   _zz_7884;
  wire       [15:0]   _zz_7885;
  wire       [31:0]   _zz_7886;
  wire       [31:0]   _zz_7887;
  wire       [15:0]   _zz_7888;
  wire       [15:0]   _zz_7889;
  wire       [15:0]   _zz_7890;
  wire       [15:0]   _zz_7891;
  wire       [15:0]   _zz_7892;
  wire       [15:0]   _zz_7893;
  wire       [15:0]   _zz_7894;
  wire       [15:0]   _zz_7895;
  wire       [15:0]   _zz_7896;
  wire       [15:0]   _zz_7897;
  wire       [15:0]   _zz_7898;
  wire       [15:0]   _zz_7899;
  wire       [15:0]   _zz_7900;
  wire       [15:0]   _zz_7901;
  wire       [15:0]   _zz_7902;
  wire       [15:0]   _zz_7903;
  wire       [15:0]   _zz_7904;
  wire       [31:0]   _zz_7905;
  wire       [31:0]   _zz_7906;
  wire       [15:0]   _zz_7907;
  wire       [31:0]   _zz_7908;
  wire       [31:0]   _zz_7909;
  wire       [15:0]   _zz_7910;
  wire       [15:0]   _zz_7911;
  wire       [15:0]   _zz_7912;
  wire       [15:0]   _zz_7913;
  wire       [15:0]   _zz_7914;
  wire       [15:0]   _zz_7915;
  wire       [15:0]   _zz_7916;
  wire       [15:0]   _zz_7917;
  wire       [15:0]   _zz_7918;
  wire       [15:0]   _zz_7919;
  wire       [15:0]   _zz_7920;
  wire       [15:0]   _zz_7921;
  wire       [15:0]   _zz_7922;
  wire       [15:0]   _zz_7923;
  wire       [15:0]   _zz_7924;
  wire       [15:0]   _zz_7925;
  wire       [15:0]   _zz_7926;
  wire       [31:0]   _zz_7927;
  wire       [31:0]   _zz_7928;
  wire       [15:0]   _zz_7929;
  wire       [31:0]   _zz_7930;
  wire       [31:0]   _zz_7931;
  wire       [15:0]   _zz_7932;
  wire       [15:0]   _zz_7933;
  wire       [15:0]   _zz_7934;
  wire       [15:0]   _zz_7935;
  wire       [15:0]   _zz_7936;
  wire       [15:0]   _zz_7937;
  wire       [15:0]   _zz_7938;
  wire       [15:0]   _zz_7939;
  wire       [15:0]   _zz_7940;
  wire       [15:0]   _zz_7941;
  wire       [15:0]   _zz_7942;
  wire       [15:0]   _zz_7943;
  wire       [15:0]   _zz_7944;
  wire       [15:0]   _zz_7945;
  wire       [15:0]   _zz_7946;
  wire       [15:0]   _zz_7947;
  wire       [15:0]   _zz_7948;
  wire       [31:0]   _zz_7949;
  wire       [31:0]   _zz_7950;
  wire       [15:0]   _zz_7951;
  wire       [31:0]   _zz_7952;
  wire       [31:0]   _zz_7953;
  wire       [15:0]   _zz_7954;
  wire       [15:0]   _zz_7955;
  wire       [15:0]   _zz_7956;
  wire       [15:0]   _zz_7957;
  wire       [15:0]   _zz_7958;
  wire       [15:0]   _zz_7959;
  wire       [15:0]   _zz_7960;
  wire       [15:0]   _zz_7961;
  wire       [15:0]   _zz_7962;
  wire       [15:0]   _zz_7963;
  wire       [15:0]   _zz_7964;
  wire       [15:0]   _zz_7965;
  wire       [15:0]   _zz_7966;
  wire       [15:0]   _zz_7967;
  wire       [15:0]   _zz_7968;
  wire       [15:0]   _zz_7969;
  wire       [15:0]   _zz_7970;
  wire       [31:0]   _zz_7971;
  wire       [31:0]   _zz_7972;
  wire       [15:0]   _zz_7973;
  wire       [31:0]   _zz_7974;
  wire       [31:0]   _zz_7975;
  wire       [15:0]   _zz_7976;
  wire       [15:0]   _zz_7977;
  wire       [15:0]   _zz_7978;
  wire       [15:0]   _zz_7979;
  wire       [15:0]   _zz_7980;
  wire       [15:0]   _zz_7981;
  wire       [15:0]   _zz_7982;
  wire       [15:0]   _zz_7983;
  wire       [15:0]   _zz_7984;
  wire       [15:0]   _zz_7985;
  wire       [15:0]   _zz_7986;
  wire       [15:0]   _zz_7987;
  wire       [15:0]   _zz_7988;
  wire       [15:0]   _zz_7989;
  wire       [15:0]   _zz_7990;
  wire       [15:0]   _zz_7991;
  wire       [15:0]   _zz_7992;
  wire       [31:0]   _zz_7993;
  wire       [31:0]   _zz_7994;
  wire       [15:0]   _zz_7995;
  wire       [31:0]   _zz_7996;
  wire       [31:0]   _zz_7997;
  wire       [15:0]   _zz_7998;
  wire       [15:0]   _zz_7999;
  wire       [15:0]   _zz_8000;
  wire       [15:0]   _zz_8001;
  wire       [15:0]   _zz_8002;
  wire       [15:0]   _zz_8003;
  wire       [15:0]   _zz_8004;
  wire       [15:0]   _zz_8005;
  wire       [15:0]   _zz_8006;
  wire       [15:0]   _zz_8007;
  wire       [15:0]   _zz_8008;
  wire       [15:0]   _zz_8009;
  wire       [15:0]   _zz_8010;
  wire       [15:0]   _zz_8011;
  wire       [15:0]   _zz_8012;
  wire       [15:0]   _zz_8013;
  wire       [15:0]   _zz_8014;
  wire       [31:0]   _zz_8015;
  wire       [31:0]   _zz_8016;
  wire       [15:0]   _zz_8017;
  wire       [31:0]   _zz_8018;
  wire       [31:0]   _zz_8019;
  wire       [15:0]   _zz_8020;
  wire       [15:0]   _zz_8021;
  wire       [15:0]   _zz_8022;
  wire       [15:0]   _zz_8023;
  wire       [15:0]   _zz_8024;
  wire       [15:0]   _zz_8025;
  wire       [15:0]   _zz_8026;
  wire       [15:0]   _zz_8027;
  wire       [15:0]   _zz_8028;
  wire       [15:0]   _zz_8029;
  wire       [15:0]   _zz_8030;
  wire       [15:0]   _zz_8031;
  wire       [15:0]   _zz_8032;
  wire       [15:0]   _zz_8033;
  wire       [15:0]   _zz_8034;
  wire       [15:0]   _zz_8035;
  wire       [15:0]   _zz_8036;
  wire       [31:0]   _zz_8037;
  wire       [31:0]   _zz_8038;
  wire       [15:0]   _zz_8039;
  wire       [31:0]   _zz_8040;
  wire       [31:0]   _zz_8041;
  wire       [15:0]   _zz_8042;
  wire       [15:0]   _zz_8043;
  wire       [15:0]   _zz_8044;
  wire       [15:0]   _zz_8045;
  wire       [15:0]   _zz_8046;
  wire       [15:0]   _zz_8047;
  wire       [15:0]   _zz_8048;
  wire       [15:0]   _zz_8049;
  wire       [15:0]   _zz_8050;
  wire       [15:0]   _zz_8051;
  wire       [15:0]   _zz_8052;
  wire       [15:0]   _zz_8053;
  wire       [15:0]   _zz_8054;
  wire       [15:0]   _zz_8055;
  wire       [15:0]   _zz_8056;
  wire       [15:0]   _zz_8057;
  wire       [15:0]   _zz_8058;
  wire       [31:0]   _zz_8059;
  wire       [31:0]   _zz_8060;
  wire       [15:0]   _zz_8061;
  wire       [31:0]   _zz_8062;
  wire       [31:0]   _zz_8063;
  wire       [15:0]   _zz_8064;
  wire       [15:0]   _zz_8065;
  wire       [15:0]   _zz_8066;
  wire       [15:0]   _zz_8067;
  wire       [15:0]   _zz_8068;
  wire       [15:0]   _zz_8069;
  wire       [15:0]   _zz_8070;
  wire       [15:0]   _zz_8071;
  wire       [15:0]   _zz_8072;
  wire       [15:0]   _zz_8073;
  wire       [15:0]   _zz_8074;
  wire       [15:0]   _zz_8075;
  wire       [15:0]   _zz_8076;
  wire       [15:0]   _zz_8077;
  wire       [15:0]   _zz_8078;
  wire       [15:0]   _zz_8079;
  wire       [15:0]   _zz_8080;
  wire       [31:0]   _zz_8081;
  wire       [31:0]   _zz_8082;
  wire       [15:0]   _zz_8083;
  wire       [31:0]   _zz_8084;
  wire       [31:0]   _zz_8085;
  wire       [15:0]   _zz_8086;
  wire       [15:0]   _zz_8087;
  wire       [15:0]   _zz_8088;
  wire       [15:0]   _zz_8089;
  wire       [15:0]   _zz_8090;
  wire       [15:0]   _zz_8091;
  wire       [15:0]   _zz_8092;
  wire       [15:0]   _zz_8093;
  wire       [15:0]   _zz_8094;
  wire       [15:0]   _zz_8095;
  wire       [15:0]   _zz_8096;
  wire       [15:0]   _zz_8097;
  wire       [15:0]   _zz_8098;
  wire       [15:0]   _zz_8099;
  wire       [15:0]   _zz_8100;
  wire       [15:0]   _zz_8101;
  wire       [15:0]   _zz_8102;
  wire       [31:0]   _zz_8103;
  wire       [31:0]   _zz_8104;
  wire       [15:0]   _zz_8105;
  wire       [31:0]   _zz_8106;
  wire       [31:0]   _zz_8107;
  wire       [15:0]   _zz_8108;
  wire       [15:0]   _zz_8109;
  wire       [15:0]   _zz_8110;
  wire       [15:0]   _zz_8111;
  wire       [15:0]   _zz_8112;
  wire       [15:0]   _zz_8113;
  wire       [15:0]   _zz_8114;
  wire       [15:0]   _zz_8115;
  wire       [15:0]   _zz_8116;
  wire       [15:0]   _zz_8117;
  wire       [15:0]   _zz_8118;
  wire       [15:0]   _zz_8119;
  wire       [15:0]   _zz_8120;
  wire       [15:0]   _zz_8121;
  wire       [15:0]   _zz_8122;
  wire       [15:0]   _zz_8123;
  wire       [15:0]   _zz_8124;
  wire       [31:0]   _zz_8125;
  wire       [31:0]   _zz_8126;
  wire       [15:0]   _zz_8127;
  wire       [31:0]   _zz_8128;
  wire       [31:0]   _zz_8129;
  wire       [15:0]   _zz_8130;
  wire       [15:0]   _zz_8131;
  wire       [15:0]   _zz_8132;
  wire       [15:0]   _zz_8133;
  wire       [15:0]   _zz_8134;
  wire       [15:0]   _zz_8135;
  wire       [15:0]   _zz_8136;
  wire       [15:0]   _zz_8137;
  wire       [15:0]   _zz_8138;
  wire       [15:0]   _zz_8139;
  wire       [15:0]   _zz_8140;
  wire       [15:0]   _zz_8141;
  wire       [15:0]   _zz_8142;
  wire       [15:0]   _zz_8143;
  wire       [15:0]   _zz_8144;
  wire       [15:0]   _zz_8145;
  wire       [15:0]   _zz_8146;
  wire       [31:0]   _zz_8147;
  wire       [31:0]   _zz_8148;
  wire       [15:0]   _zz_8149;
  wire       [31:0]   _zz_8150;
  wire       [31:0]   _zz_8151;
  wire       [15:0]   _zz_8152;
  wire       [15:0]   _zz_8153;
  wire       [15:0]   _zz_8154;
  wire       [15:0]   _zz_8155;
  wire       [15:0]   _zz_8156;
  wire       [15:0]   _zz_8157;
  wire       [15:0]   _zz_8158;
  wire       [15:0]   _zz_8159;
  wire       [15:0]   _zz_8160;
  wire       [15:0]   _zz_8161;
  wire       [15:0]   _zz_8162;
  wire       [15:0]   _zz_8163;
  wire       [15:0]   _zz_8164;
  wire       [15:0]   _zz_8165;
  wire       [15:0]   _zz_8166;
  wire       [15:0]   _zz_8167;
  wire       [15:0]   _zz_8168;
  wire       [31:0]   _zz_8169;
  wire       [31:0]   _zz_8170;
  wire       [15:0]   _zz_8171;
  wire       [31:0]   _zz_8172;
  wire       [31:0]   _zz_8173;
  wire       [15:0]   _zz_8174;
  wire       [15:0]   _zz_8175;
  wire       [15:0]   _zz_8176;
  wire       [15:0]   _zz_8177;
  wire       [15:0]   _zz_8178;
  wire       [15:0]   _zz_8179;
  wire       [15:0]   _zz_8180;
  wire       [15:0]   _zz_8181;
  wire       [15:0]   _zz_8182;
  wire       [15:0]   _zz_8183;
  wire       [15:0]   _zz_8184;
  wire       [15:0]   _zz_8185;
  wire       [15:0]   _zz_8186;
  wire       [15:0]   _zz_8187;
  wire       [15:0]   _zz_8188;
  wire       [15:0]   _zz_8189;
  wire       [15:0]   _zz_8190;
  wire       [31:0]   _zz_8191;
  wire       [31:0]   _zz_8192;
  wire       [15:0]   _zz_8193;
  wire       [31:0]   _zz_8194;
  wire       [31:0]   _zz_8195;
  wire       [15:0]   _zz_8196;
  wire       [15:0]   _zz_8197;
  wire       [15:0]   _zz_8198;
  wire       [15:0]   _zz_8199;
  wire       [15:0]   _zz_8200;
  wire       [15:0]   _zz_8201;
  wire       [15:0]   _zz_8202;
  wire       [15:0]   _zz_8203;
  wire       [15:0]   _zz_8204;
  wire       [15:0]   _zz_8205;
  wire       [15:0]   _zz_8206;
  wire       [15:0]   _zz_8207;
  wire       [15:0]   _zz_8208;
  wire       [15:0]   _zz_8209;
  wire       [15:0]   _zz_8210;
  wire       [15:0]   _zz_8211;
  wire       [15:0]   _zz_8212;
  wire       [31:0]   _zz_8213;
  wire       [31:0]   _zz_8214;
  wire       [15:0]   _zz_8215;
  wire       [31:0]   _zz_8216;
  wire       [31:0]   _zz_8217;
  wire       [15:0]   _zz_8218;
  wire       [15:0]   _zz_8219;
  wire       [15:0]   _zz_8220;
  wire       [15:0]   _zz_8221;
  wire       [15:0]   _zz_8222;
  wire       [15:0]   _zz_8223;
  wire       [15:0]   _zz_8224;
  wire       [15:0]   _zz_8225;
  wire       [15:0]   _zz_8226;
  wire       [15:0]   _zz_8227;
  wire       [15:0]   _zz_8228;
  wire       [15:0]   _zz_8229;
  wire       [15:0]   _zz_8230;
  wire       [15:0]   _zz_8231;
  wire       [15:0]   _zz_8232;
  wire       [15:0]   _zz_8233;
  wire       [15:0]   _zz_8234;
  wire       [31:0]   _zz_8235;
  wire       [31:0]   _zz_8236;
  wire       [15:0]   _zz_8237;
  wire       [31:0]   _zz_8238;
  wire       [31:0]   _zz_8239;
  wire       [15:0]   _zz_8240;
  wire       [15:0]   _zz_8241;
  wire       [15:0]   _zz_8242;
  wire       [15:0]   _zz_8243;
  wire       [15:0]   _zz_8244;
  wire       [15:0]   _zz_8245;
  wire       [15:0]   _zz_8246;
  wire       [15:0]   _zz_8247;
  wire       [15:0]   _zz_8248;
  wire       [15:0]   _zz_8249;
  wire       [15:0]   _zz_8250;
  wire       [15:0]   _zz_8251;
  wire       [15:0]   _zz_8252;
  wire       [15:0]   _zz_8253;
  wire       [15:0]   _zz_8254;
  wire       [15:0]   _zz_8255;
  wire       [15:0]   _zz_8256;
  wire       [31:0]   _zz_8257;
  wire       [31:0]   _zz_8258;
  wire       [15:0]   _zz_8259;
  wire       [31:0]   _zz_8260;
  wire       [31:0]   _zz_8261;
  wire       [15:0]   _zz_8262;
  wire       [15:0]   _zz_8263;
  wire       [15:0]   _zz_8264;
  wire       [15:0]   _zz_8265;
  wire       [15:0]   _zz_8266;
  wire       [15:0]   _zz_8267;
  wire       [15:0]   _zz_8268;
  wire       [15:0]   _zz_8269;
  wire       [15:0]   _zz_8270;
  wire       [15:0]   _zz_8271;
  wire       [15:0]   _zz_8272;
  wire       [15:0]   _zz_8273;
  wire       [15:0]   _zz_8274;
  wire       [15:0]   _zz_8275;
  wire       [15:0]   _zz_8276;
  wire       [15:0]   _zz_8277;
  wire       [15:0]   _zz_8278;
  wire       [31:0]   _zz_8279;
  wire       [31:0]   _zz_8280;
  wire       [15:0]   _zz_8281;
  wire       [31:0]   _zz_8282;
  wire       [31:0]   _zz_8283;
  wire       [15:0]   _zz_8284;
  wire       [15:0]   _zz_8285;
  wire       [15:0]   _zz_8286;
  wire       [15:0]   _zz_8287;
  wire       [15:0]   _zz_8288;
  wire       [15:0]   _zz_8289;
  wire       [15:0]   _zz_8290;
  wire       [15:0]   _zz_8291;
  wire       [15:0]   _zz_8292;
  wire       [15:0]   _zz_8293;
  wire       [15:0]   _zz_8294;
  wire       [15:0]   _zz_8295;
  wire       [15:0]   _zz_8296;
  wire       [15:0]   _zz_8297;
  wire       [15:0]   _zz_8298;
  wire       [15:0]   _zz_8299;
  wire       [15:0]   _zz_8300;
  wire       [31:0]   _zz_8301;
  wire       [31:0]   _zz_8302;
  wire       [15:0]   _zz_8303;
  wire       [31:0]   _zz_8304;
  wire       [31:0]   _zz_8305;
  wire       [15:0]   _zz_8306;
  wire       [15:0]   _zz_8307;
  wire       [15:0]   _zz_8308;
  wire       [15:0]   _zz_8309;
  wire       [15:0]   _zz_8310;
  wire       [15:0]   _zz_8311;
  wire       [15:0]   _zz_8312;
  wire       [15:0]   _zz_8313;
  wire       [15:0]   _zz_8314;
  wire       [15:0]   _zz_8315;
  wire       [15:0]   _zz_8316;
  wire       [15:0]   _zz_8317;
  wire       [15:0]   _zz_8318;
  wire       [15:0]   _zz_8319;
  wire       [15:0]   _zz_8320;
  wire       [15:0]   _zz_8321;
  wire       [15:0]   _zz_8322;
  wire       [31:0]   _zz_8323;
  wire       [31:0]   _zz_8324;
  wire       [15:0]   _zz_8325;
  wire       [31:0]   _zz_8326;
  wire       [31:0]   _zz_8327;
  wire       [15:0]   _zz_8328;
  wire       [15:0]   _zz_8329;
  wire       [15:0]   _zz_8330;
  wire       [15:0]   _zz_8331;
  wire       [15:0]   _zz_8332;
  wire       [15:0]   _zz_8333;
  wire       [15:0]   _zz_8334;
  wire       [15:0]   _zz_8335;
  wire       [15:0]   _zz_8336;
  wire       [15:0]   _zz_8337;
  wire       [15:0]   _zz_8338;
  wire       [15:0]   _zz_8339;
  wire       [15:0]   _zz_8340;
  wire       [15:0]   _zz_8341;
  wire       [15:0]   _zz_8342;
  wire       [15:0]   _zz_8343;
  wire       [15:0]   _zz_8344;
  wire       [31:0]   _zz_8345;
  wire       [31:0]   _zz_8346;
  wire       [15:0]   _zz_8347;
  wire       [31:0]   _zz_8348;
  wire       [31:0]   _zz_8349;
  wire       [15:0]   _zz_8350;
  wire       [15:0]   _zz_8351;
  wire       [15:0]   _zz_8352;
  wire       [15:0]   _zz_8353;
  wire       [15:0]   _zz_8354;
  wire       [15:0]   _zz_8355;
  wire       [15:0]   _zz_8356;
  wire       [15:0]   _zz_8357;
  wire       [15:0]   _zz_8358;
  wire       [15:0]   _zz_8359;
  wire       [15:0]   _zz_8360;
  wire       [15:0]   _zz_8361;
  wire       [15:0]   _zz_8362;
  wire       [15:0]   _zz_8363;
  wire       [15:0]   _zz_8364;
  wire       [15:0]   _zz_8365;
  wire       [15:0]   _zz_8366;
  wire       [31:0]   _zz_8367;
  wire       [31:0]   _zz_8368;
  wire       [15:0]   _zz_8369;
  wire       [31:0]   _zz_8370;
  wire       [31:0]   _zz_8371;
  wire       [15:0]   _zz_8372;
  wire       [15:0]   _zz_8373;
  wire       [15:0]   _zz_8374;
  wire       [15:0]   _zz_8375;
  wire       [15:0]   _zz_8376;
  wire       [15:0]   _zz_8377;
  wire       [15:0]   _zz_8378;
  wire       [15:0]   _zz_8379;
  wire       [15:0]   _zz_8380;
  wire       [15:0]   _zz_8381;
  wire       [15:0]   _zz_8382;
  wire       [15:0]   _zz_8383;
  wire       [15:0]   _zz_8384;
  wire       [15:0]   _zz_8385;
  wire       [15:0]   _zz_8386;
  wire       [15:0]   _zz_8387;
  wire       [15:0]   _zz_8388;
  wire       [31:0]   _zz_8389;
  wire       [31:0]   _zz_8390;
  wire       [15:0]   _zz_8391;
  wire       [31:0]   _zz_8392;
  wire       [31:0]   _zz_8393;
  wire       [15:0]   _zz_8394;
  wire       [15:0]   _zz_8395;
  wire       [15:0]   _zz_8396;
  wire       [15:0]   _zz_8397;
  wire       [15:0]   _zz_8398;
  wire       [15:0]   _zz_8399;
  wire       [15:0]   _zz_8400;
  wire       [15:0]   _zz_8401;
  wire       [15:0]   _zz_8402;
  wire       [15:0]   _zz_8403;
  wire       [15:0]   _zz_8404;
  wire       [15:0]   _zz_8405;
  wire       [15:0]   _zz_8406;
  wire       [15:0]   _zz_8407;
  wire       [15:0]   _zz_8408;
  wire       [15:0]   _zz_8409;
  wire       [15:0]   _zz_8410;
  wire       [31:0]   _zz_8411;
  wire       [31:0]   _zz_8412;
  wire       [15:0]   _zz_8413;
  wire       [31:0]   _zz_8414;
  wire       [31:0]   _zz_8415;
  wire       [15:0]   _zz_8416;
  wire       [15:0]   _zz_8417;
  wire       [15:0]   _zz_8418;
  wire       [15:0]   _zz_8419;
  wire       [15:0]   _zz_8420;
  wire       [15:0]   _zz_8421;
  wire       [15:0]   _zz_8422;
  wire       [15:0]   _zz_8423;
  wire       [15:0]   _zz_8424;
  wire       [15:0]   _zz_8425;
  wire       [15:0]   _zz_8426;
  wire       [15:0]   _zz_8427;
  wire       [15:0]   _zz_8428;
  wire       [15:0]   _zz_8429;
  wire       [15:0]   _zz_8430;
  wire       [15:0]   _zz_8431;
  wire       [15:0]   _zz_8432;
  wire       [31:0]   _zz_8433;
  wire       [31:0]   _zz_8434;
  wire       [15:0]   _zz_8435;
  wire       [31:0]   _zz_8436;
  wire       [31:0]   _zz_8437;
  wire       [15:0]   _zz_8438;
  wire       [15:0]   _zz_8439;
  wire       [15:0]   _zz_8440;
  wire       [15:0]   _zz_8441;
  wire       [15:0]   _zz_8442;
  wire       [15:0]   _zz_8443;
  wire       [15:0]   _zz_8444;
  wire       [15:0]   _zz_8445;
  wire       [15:0]   _zz_8446;
  wire       [15:0]   _zz_8447;
  wire       [15:0]   _zz_8448;
  wire       [15:0]   _zz_8449;
  wire       [15:0]   _zz_8450;
  wire       [15:0]   _zz_8451;
  wire       [15:0]   _zz_8452;
  wire       [15:0]   _zz_8453;
  wire       [15:0]   _zz_8454;
  wire       [31:0]   _zz_8455;
  wire       [31:0]   _zz_8456;
  wire       [15:0]   _zz_8457;
  wire       [31:0]   _zz_8458;
  wire       [31:0]   _zz_8459;
  wire       [15:0]   _zz_8460;
  wire       [15:0]   _zz_8461;
  wire       [15:0]   _zz_8462;
  wire       [15:0]   _zz_8463;
  wire       [15:0]   _zz_8464;
  wire       [15:0]   _zz_8465;
  wire       [15:0]   _zz_8466;
  wire       [15:0]   _zz_8467;
  wire       [15:0]   _zz_8468;
  wire       [15:0]   _zz_8469;
  wire       [15:0]   _zz_8470;
  wire       [15:0]   _zz_8471;
  wire       [15:0]   _zz_8472;
  wire       [15:0]   _zz_8473;
  wire       [15:0]   _zz_8474;
  wire       [15:0]   _zz_8475;
  wire       [15:0]   _zz_8476;
  wire       [31:0]   _zz_8477;
  wire       [31:0]   _zz_8478;
  wire       [15:0]   _zz_8479;
  wire       [31:0]   _zz_8480;
  wire       [31:0]   _zz_8481;
  wire       [15:0]   _zz_8482;
  wire       [15:0]   _zz_8483;
  wire       [15:0]   _zz_8484;
  wire       [15:0]   _zz_8485;
  wire       [15:0]   _zz_8486;
  wire       [15:0]   _zz_8487;
  wire       [15:0]   _zz_8488;
  wire       [15:0]   _zz_8489;
  wire       [15:0]   _zz_8490;
  wire       [15:0]   _zz_8491;
  wire       [15:0]   _zz_8492;
  wire       [15:0]   _zz_8493;
  wire       [15:0]   _zz_8494;
  wire       [15:0]   _zz_8495;
  wire       [15:0]   _zz_8496;
  wire       [15:0]   _zz_8497;
  wire       [15:0]   _zz_8498;
  wire       [31:0]   _zz_8499;
  wire       [31:0]   _zz_8500;
  wire       [15:0]   _zz_8501;
  wire       [31:0]   _zz_8502;
  wire       [31:0]   _zz_8503;
  wire       [15:0]   _zz_8504;
  wire       [15:0]   _zz_8505;
  wire       [15:0]   _zz_8506;
  wire       [15:0]   _zz_8507;
  wire       [15:0]   _zz_8508;
  wire       [15:0]   _zz_8509;
  wire       [15:0]   _zz_8510;
  wire       [15:0]   _zz_8511;
  wire       [15:0]   _zz_8512;
  wire       [15:0]   _zz_8513;
  wire       [15:0]   _zz_8514;
  wire       [15:0]   _zz_8515;
  wire       [15:0]   _zz_8516;
  wire       [15:0]   _zz_8517;
  wire       [15:0]   _zz_8518;
  wire       [15:0]   _zz_8519;
  wire       [15:0]   _zz_8520;
  wire       [31:0]   _zz_8521;
  wire       [31:0]   _zz_8522;
  wire       [15:0]   _zz_8523;
  wire       [31:0]   _zz_8524;
  wire       [31:0]   _zz_8525;
  wire       [15:0]   _zz_8526;
  wire       [15:0]   _zz_8527;
  wire       [15:0]   _zz_8528;
  wire       [15:0]   _zz_8529;
  wire       [15:0]   _zz_8530;
  wire       [15:0]   _zz_8531;
  wire       [15:0]   _zz_8532;
  wire       [15:0]   _zz_8533;
  wire       [15:0]   _zz_8534;
  wire       [15:0]   _zz_8535;
  wire       [15:0]   _zz_8536;
  wire       [15:0]   _zz_8537;
  wire       [15:0]   _zz_8538;
  wire       [15:0]   _zz_8539;
  wire       [15:0]   _zz_8540;
  wire       [15:0]   _zz_8541;
  wire       [15:0]   _zz_8542;
  wire       [31:0]   _zz_8543;
  wire       [31:0]   _zz_8544;
  wire       [15:0]   _zz_8545;
  wire       [31:0]   _zz_8546;
  wire       [31:0]   _zz_8547;
  wire       [15:0]   _zz_8548;
  wire       [15:0]   _zz_8549;
  wire       [15:0]   _zz_8550;
  wire       [15:0]   _zz_8551;
  wire       [15:0]   _zz_8552;
  wire       [15:0]   _zz_8553;
  wire       [15:0]   _zz_8554;
  wire       [15:0]   _zz_8555;
  wire       [15:0]   _zz_8556;
  wire       [15:0]   _zz_8557;
  wire       [15:0]   _zz_8558;
  wire       [15:0]   _zz_8559;
  wire       [15:0]   _zz_8560;
  wire       [15:0]   _zz_8561;
  wire       [15:0]   _zz_8562;
  wire       [15:0]   _zz_8563;
  wire       [15:0]   _zz_8564;
  wire       [31:0]   _zz_8565;
  wire       [31:0]   _zz_8566;
  wire       [15:0]   _zz_8567;
  wire       [31:0]   _zz_8568;
  wire       [31:0]   _zz_8569;
  wire       [15:0]   _zz_8570;
  wire       [15:0]   _zz_8571;
  wire       [15:0]   _zz_8572;
  wire       [15:0]   _zz_8573;
  wire       [15:0]   _zz_8574;
  wire       [15:0]   _zz_8575;
  wire       [15:0]   _zz_8576;
  wire       [15:0]   _zz_8577;
  wire       [15:0]   _zz_8578;
  wire       [15:0]   _zz_8579;
  wire       [15:0]   _zz_8580;
  wire       [15:0]   _zz_8581;
  wire       [15:0]   _zz_8582;
  wire       [15:0]   _zz_8583;
  wire       [15:0]   _zz_8584;
  wire       [15:0]   _zz_8585;
  wire       [15:0]   _zz_8586;
  wire       [31:0]   _zz_8587;
  wire       [31:0]   _zz_8588;
  wire       [15:0]   _zz_8589;
  wire       [31:0]   _zz_8590;
  wire       [31:0]   _zz_8591;
  wire       [15:0]   _zz_8592;
  wire       [15:0]   _zz_8593;
  wire       [15:0]   _zz_8594;
  wire       [15:0]   _zz_8595;
  wire       [15:0]   _zz_8596;
  wire       [15:0]   _zz_8597;
  wire       [15:0]   _zz_8598;
  wire       [15:0]   _zz_8599;
  wire       [15:0]   _zz_8600;
  wire       [15:0]   _zz_8601;
  wire       [15:0]   _zz_8602;
  wire       [15:0]   _zz_8603;
  wire       [15:0]   _zz_8604;
  wire       [15:0]   _zz_8605;
  wire       [15:0]   _zz_8606;
  wire       [15:0]   _zz_8607;
  wire       [15:0]   _zz_8608;
  wire       [31:0]   _zz_8609;
  wire       [31:0]   _zz_8610;
  wire       [15:0]   _zz_8611;
  wire       [31:0]   _zz_8612;
  wire       [31:0]   _zz_8613;
  wire       [15:0]   _zz_8614;
  wire       [15:0]   _zz_8615;
  wire       [15:0]   _zz_8616;
  wire       [15:0]   _zz_8617;
  wire       [15:0]   _zz_8618;
  wire       [15:0]   _zz_8619;
  wire       [15:0]   _zz_8620;
  wire       [15:0]   _zz_8621;
  wire       [15:0]   _zz_8622;
  wire       [15:0]   _zz_8623;
  wire       [15:0]   _zz_8624;
  wire       [15:0]   _zz_8625;
  wire       [15:0]   _zz_8626;
  wire       [15:0]   _zz_8627;
  wire       [15:0]   _zz_8628;
  wire       [15:0]   _zz_8629;
  wire       [15:0]   _zz_8630;
  wire       [31:0]   _zz_8631;
  wire       [31:0]   _zz_8632;
  wire       [15:0]   _zz_8633;
  wire       [31:0]   _zz_8634;
  wire       [31:0]   _zz_8635;
  wire       [15:0]   _zz_8636;
  wire       [15:0]   _zz_8637;
  wire       [15:0]   _zz_8638;
  wire       [15:0]   _zz_8639;
  wire       [15:0]   _zz_8640;
  wire       [15:0]   _zz_8641;
  wire       [15:0]   _zz_8642;
  wire       [15:0]   _zz_8643;
  wire       [15:0]   _zz_8644;
  wire       [15:0]   _zz_8645;
  wire       [15:0]   _zz_8646;
  wire       [15:0]   _zz_8647;
  wire       [15:0]   _zz_8648;
  wire       [15:0]   _zz_8649;
  wire       [15:0]   _zz_8650;
  wire       [15:0]   _zz_8651;
  wire       [15:0]   _zz_8652;
  wire       [31:0]   _zz_8653;
  wire       [31:0]   _zz_8654;
  wire       [15:0]   _zz_8655;
  wire       [31:0]   _zz_8656;
  wire       [31:0]   _zz_8657;
  wire       [15:0]   _zz_8658;
  wire       [15:0]   _zz_8659;
  wire       [15:0]   _zz_8660;
  wire       [15:0]   _zz_8661;
  wire       [15:0]   _zz_8662;
  wire       [15:0]   _zz_8663;
  wire       [15:0]   _zz_8664;
  wire       [15:0]   _zz_8665;
  wire       [15:0]   _zz_8666;
  wire       [15:0]   _zz_8667;
  wire       [15:0]   _zz_8668;
  wire       [15:0]   _zz_8669;
  wire       [15:0]   _zz_8670;
  wire       [15:0]   _zz_8671;
  wire       [15:0]   _zz_8672;
  wire       [15:0]   _zz_8673;
  wire       [15:0]   _zz_8674;
  wire       [31:0]   _zz_8675;
  wire       [31:0]   _zz_8676;
  wire       [15:0]   _zz_8677;
  wire       [31:0]   _zz_8678;
  wire       [31:0]   _zz_8679;
  wire       [15:0]   _zz_8680;
  wire       [15:0]   _zz_8681;
  wire       [15:0]   _zz_8682;
  wire       [15:0]   _zz_8683;
  wire       [15:0]   _zz_8684;
  wire       [15:0]   _zz_8685;
  wire       [15:0]   _zz_8686;
  wire       [15:0]   _zz_8687;
  wire       [15:0]   _zz_8688;
  wire       [15:0]   _zz_8689;
  wire       [15:0]   _zz_8690;
  wire       [15:0]   _zz_8691;
  wire       [15:0]   _zz_8692;
  wire       [15:0]   _zz_8693;
  wire       [15:0]   _zz_8694;
  wire       [15:0]   _zz_8695;
  wire       [15:0]   _zz_8696;
  wire       [31:0]   _zz_8697;
  wire       [31:0]   _zz_8698;
  wire       [15:0]   _zz_8699;
  wire       [31:0]   _zz_8700;
  wire       [31:0]   _zz_8701;
  wire       [15:0]   _zz_8702;
  wire       [15:0]   _zz_8703;
  wire       [15:0]   _zz_8704;
  wire       [15:0]   _zz_8705;
  wire       [15:0]   _zz_8706;
  wire       [15:0]   _zz_8707;
  wire       [15:0]   _zz_8708;
  wire       [15:0]   _zz_8709;
  wire       [15:0]   _zz_8710;
  wire       [15:0]   _zz_8711;
  wire       [15:0]   _zz_8712;
  wire       [15:0]   _zz_8713;
  wire       [15:0]   _zz_8714;
  wire       [15:0]   _zz_8715;
  wire       [15:0]   _zz_8716;
  wire       [15:0]   _zz_8717;
  wire       [15:0]   _zz_8718;
  wire       [31:0]   _zz_8719;
  wire       [31:0]   _zz_8720;
  wire       [15:0]   _zz_8721;
  wire       [31:0]   _zz_8722;
  wire       [31:0]   _zz_8723;
  wire       [15:0]   _zz_8724;
  wire       [15:0]   _zz_8725;
  wire       [15:0]   _zz_8726;
  wire       [15:0]   _zz_8727;
  wire       [15:0]   _zz_8728;
  wire       [15:0]   _zz_8729;
  wire       [15:0]   _zz_8730;
  wire       [15:0]   _zz_8731;
  wire       [15:0]   _zz_8732;
  wire       [15:0]   _zz_8733;
  wire       [15:0]   _zz_8734;
  wire       [15:0]   _zz_8735;
  wire       [15:0]   _zz_8736;
  wire       [15:0]   _zz_8737;
  wire       [15:0]   _zz_8738;
  wire       [15:0]   _zz_8739;
  wire       [15:0]   _zz_8740;
  wire       [31:0]   _zz_8741;
  wire       [31:0]   _zz_8742;
  wire       [15:0]   _zz_8743;
  wire       [31:0]   _zz_8744;
  wire       [31:0]   _zz_8745;
  wire       [15:0]   _zz_8746;
  wire       [15:0]   _zz_8747;
  wire       [15:0]   _zz_8748;
  wire       [15:0]   _zz_8749;
  wire       [15:0]   _zz_8750;
  wire       [15:0]   _zz_8751;
  wire       [15:0]   _zz_8752;
  wire       [15:0]   _zz_8753;
  wire       [15:0]   _zz_8754;
  wire       [15:0]   _zz_8755;
  wire       [15:0]   _zz_8756;
  wire       [15:0]   _zz_8757;
  wire       [15:0]   _zz_8758;
  wire       [15:0]   _zz_8759;
  wire       [15:0]   _zz_8760;
  wire       [15:0]   _zz_8761;
  wire       [15:0]   _zz_8762;
  wire       [31:0]   _zz_8763;
  wire       [31:0]   _zz_8764;
  wire       [15:0]   _zz_8765;
  wire       [31:0]   _zz_8766;
  wire       [31:0]   _zz_8767;
  wire       [15:0]   _zz_8768;
  wire       [15:0]   _zz_8769;
  wire       [15:0]   _zz_8770;
  wire       [15:0]   _zz_8771;
  wire       [15:0]   _zz_8772;
  wire       [15:0]   _zz_8773;
  wire       [15:0]   _zz_8774;
  wire       [15:0]   _zz_8775;
  wire       [15:0]   _zz_8776;
  wire       [15:0]   _zz_8777;
  wire       [15:0]   _zz_8778;
  wire       [15:0]   _zz_8779;
  wire       [15:0]   _zz_8780;
  wire       [15:0]   _zz_8781;
  wire       [15:0]   _zz_8782;
  wire       [15:0]   _zz_8783;
  wire       [15:0]   _zz_8784;
  wire       [31:0]   _zz_8785;
  wire       [31:0]   _zz_8786;
  wire       [15:0]   _zz_8787;
  wire       [31:0]   _zz_8788;
  wire       [31:0]   _zz_8789;
  wire       [15:0]   _zz_8790;
  wire       [15:0]   _zz_8791;
  wire       [15:0]   _zz_8792;
  wire       [15:0]   _zz_8793;
  wire       [15:0]   _zz_8794;
  wire       [15:0]   _zz_8795;
  wire       [15:0]   _zz_8796;
  wire       [15:0]   _zz_8797;
  wire       [15:0]   _zz_8798;
  wire       [15:0]   _zz_8799;
  wire       [15:0]   _zz_8800;
  wire       [15:0]   _zz_8801;
  wire       [15:0]   _zz_8802;
  wire       [15:0]   _zz_8803;
  wire       [15:0]   _zz_8804;
  wire       [15:0]   _zz_8805;
  wire       [15:0]   _zz_8806;
  wire       [31:0]   _zz_8807;
  wire       [31:0]   _zz_8808;
  wire       [15:0]   _zz_8809;
  wire       [31:0]   _zz_8810;
  wire       [31:0]   _zz_8811;
  wire       [15:0]   _zz_8812;
  wire       [15:0]   _zz_8813;
  wire       [15:0]   _zz_8814;
  wire       [15:0]   _zz_8815;
  wire       [15:0]   _zz_8816;
  wire       [15:0]   _zz_8817;
  wire       [15:0]   _zz_8818;
  wire       [15:0]   _zz_8819;
  wire       [15:0]   _zz_8820;
  wire       [15:0]   _zz_8821;
  wire       [15:0]   _zz_8822;
  wire       [15:0]   _zz_8823;
  wire       [15:0]   _zz_8824;
  wire       [15:0]   _zz_8825;
  wire       [15:0]   _zz_8826;
  wire       [15:0]   _zz_8827;
  wire       [15:0]   _zz_8828;
  wire       [31:0]   _zz_8829;
  wire       [31:0]   _zz_8830;
  wire       [15:0]   _zz_8831;
  wire       [31:0]   _zz_8832;
  wire       [31:0]   _zz_8833;
  wire       [15:0]   _zz_8834;
  wire       [15:0]   _zz_8835;
  wire       [15:0]   _zz_8836;
  wire       [15:0]   _zz_8837;
  wire       [15:0]   _zz_8838;
  wire       [15:0]   _zz_8839;
  wire       [15:0]   _zz_8840;
  wire       [15:0]   _zz_8841;
  wire       [15:0]   _zz_8842;
  wire       [15:0]   _zz_8843;
  wire       [15:0]   _zz_8844;
  wire       [15:0]   _zz_8845;
  wire       [15:0]   _zz_8846;
  wire       [15:0]   _zz_8847;
  wire       [15:0]   _zz_8848;
  wire       [15:0]   _zz_8849;
  wire       [15:0]   _zz_8850;
  wire       [31:0]   _zz_8851;
  wire       [31:0]   _zz_8852;
  wire       [15:0]   _zz_8853;
  wire       [31:0]   _zz_8854;
  wire       [31:0]   _zz_8855;
  wire       [15:0]   _zz_8856;
  wire       [15:0]   _zz_8857;
  wire       [15:0]   _zz_8858;
  wire       [15:0]   _zz_8859;
  wire       [15:0]   _zz_8860;
  wire       [15:0]   _zz_8861;
  wire       [15:0]   _zz_8862;
  wire       [15:0]   _zz_8863;
  wire       [15:0]   _zz_8864;
  wire       [15:0]   _zz_8865;
  wire       [15:0]   _zz_8866;
  wire       [15:0]   _zz_8867;
  wire       [15:0]   _zz_8868;
  wire       [15:0]   _zz_8869;
  wire       [15:0]   _zz_8870;
  wire       [15:0]   _zz_8871;
  wire       [15:0]   _zz_8872;
  wire       [31:0]   _zz_8873;
  wire       [31:0]   _zz_8874;
  wire       [15:0]   _zz_8875;
  wire       [31:0]   _zz_8876;
  wire       [31:0]   _zz_8877;
  wire       [15:0]   _zz_8878;
  wire       [15:0]   _zz_8879;
  wire       [15:0]   _zz_8880;
  wire       [15:0]   _zz_8881;
  wire       [15:0]   _zz_8882;
  wire       [15:0]   _zz_8883;
  wire       [15:0]   _zz_8884;
  wire       [15:0]   _zz_8885;
  wire       [15:0]   _zz_8886;
  wire       [15:0]   _zz_8887;
  wire       [15:0]   _zz_8888;
  wire       [15:0]   _zz_8889;
  wire       [15:0]   _zz_8890;
  wire       [15:0]   _zz_8891;
  wire       [15:0]   _zz_8892;
  wire       [15:0]   _zz_8893;
  wire       [15:0]   _zz_8894;
  wire       [31:0]   _zz_8895;
  wire       [31:0]   _zz_8896;
  wire       [15:0]   _zz_8897;
  wire       [31:0]   _zz_8898;
  wire       [31:0]   _zz_8899;
  wire       [15:0]   _zz_8900;
  wire       [15:0]   _zz_8901;
  wire       [15:0]   _zz_8902;
  wire       [15:0]   _zz_8903;
  wire       [15:0]   _zz_8904;
  wire       [15:0]   _zz_8905;
  wire       [15:0]   _zz_8906;
  wire       [15:0]   _zz_8907;
  wire       [15:0]   _zz_8908;
  wire       [15:0]   _zz_8909;
  wire       [15:0]   _zz_8910;
  wire       [15:0]   _zz_8911;
  wire       [15:0]   _zz_8912;
  wire       [15:0]   _zz_8913;
  wire       [15:0]   _zz_8914;
  wire       [15:0]   _zz_8915;
  wire       [15:0]   _zz_8916;
  wire       [31:0]   _zz_8917;
  wire       [31:0]   _zz_8918;
  wire       [15:0]   _zz_8919;
  wire       [31:0]   _zz_8920;
  wire       [31:0]   _zz_8921;
  wire       [15:0]   _zz_8922;
  wire       [15:0]   _zz_8923;
  wire       [15:0]   _zz_8924;
  wire       [15:0]   _zz_8925;
  wire       [15:0]   _zz_8926;
  wire       [15:0]   _zz_8927;
  wire       [15:0]   _zz_8928;
  wire       [15:0]   _zz_8929;
  wire       [15:0]   _zz_8930;
  wire       [15:0]   _zz_8931;
  wire       [15:0]   _zz_8932;
  wire       [15:0]   _zz_8933;
  wire       [15:0]   _zz_8934;
  wire       [15:0]   _zz_8935;
  wire       [15:0]   _zz_8936;
  wire       [15:0]   _zz_8937;
  wire       [15:0]   _zz_8938;
  wire       [31:0]   _zz_8939;
  wire       [31:0]   _zz_8940;
  wire       [15:0]   _zz_8941;
  wire       [31:0]   _zz_8942;
  wire       [31:0]   _zz_8943;
  wire       [15:0]   _zz_8944;
  wire       [15:0]   _zz_8945;
  wire       [15:0]   _zz_8946;
  wire       [15:0]   _zz_8947;
  wire       [15:0]   _zz_8948;
  wire       [15:0]   _zz_8949;
  wire       [15:0]   _zz_8950;
  wire       [15:0]   _zz_8951;
  wire       [15:0]   _zz_8952;
  wire       [15:0]   _zz_8953;
  wire       [15:0]   _zz_8954;
  wire       [15:0]   _zz_8955;
  wire       [15:0]   _zz_8956;
  wire       [15:0]   _zz_8957;
  wire       [15:0]   _zz_8958;
  wire       [15:0]   _zz_8959;
  wire       [15:0]   _zz_8960;
  wire       [31:0]   _zz_8961;
  wire       [31:0]   _zz_8962;
  wire       [15:0]   _zz_8963;
  wire       [31:0]   _zz_8964;
  wire       [31:0]   _zz_8965;
  wire       [15:0]   _zz_8966;
  wire       [15:0]   _zz_8967;
  wire       [15:0]   _zz_8968;
  wire       [15:0]   _zz_8969;
  wire       [15:0]   _zz_8970;
  wire       [15:0]   _zz_8971;
  wire       [15:0]   _zz_8972;
  wire       [15:0]   _zz_8973;
  wire       [15:0]   _zz_8974;
  wire       [15:0]   _zz_8975;
  wire       [15:0]   _zz_8976;
  wire       [15:0]   _zz_8977;
  wire       [15:0]   _zz_8978;
  wire       [15:0]   _zz_8979;
  wire       [15:0]   _zz_8980;
  wire       [15:0]   _zz_8981;
  wire       [15:0]   _zz_8982;
  wire       [31:0]   _zz_8983;
  wire       [31:0]   _zz_8984;
  wire       [15:0]   _zz_8985;
  wire       [31:0]   _zz_8986;
  wire       [31:0]   _zz_8987;
  wire       [15:0]   _zz_8988;
  wire       [15:0]   _zz_8989;
  wire       [15:0]   _zz_8990;
  wire       [15:0]   _zz_8991;
  wire       [15:0]   _zz_8992;
  wire       [15:0]   _zz_8993;
  wire       [15:0]   _zz_8994;
  wire       [15:0]   _zz_8995;
  wire       [15:0]   _zz_8996;
  wire       [15:0]   _zz_8997;
  wire       [15:0]   _zz_8998;
  wire       [15:0]   _zz_8999;
  wire       [15:0]   _zz_9000;
  wire       [15:0]   _zz_9001;
  wire       [15:0]   _zz_9002;
  wire       [15:0]   _zz_9003;
  wire       [15:0]   _zz_9004;
  wire       [31:0]   _zz_9005;
  wire       [31:0]   _zz_9006;
  wire       [15:0]   _zz_9007;
  wire       [31:0]   _zz_9008;
  wire       [31:0]   _zz_9009;
  wire       [15:0]   _zz_9010;
  wire       [15:0]   _zz_9011;
  wire       [15:0]   _zz_9012;
  wire       [15:0]   _zz_9013;
  wire       [15:0]   _zz_9014;
  wire       [15:0]   _zz_9015;
  wire       [15:0]   _zz_9016;
  wire       [15:0]   _zz_9017;
  wire       [15:0]   _zz_9018;
  wire       [15:0]   _zz_9019;
  wire       [15:0]   _zz_9020;
  wire       [15:0]   _zz_9021;
  wire       [15:0]   _zz_9022;
  wire       [15:0]   _zz_9023;
  wire       [15:0]   _zz_9024;
  wire       [15:0]   _zz_9025;
  wire       [15:0]   _zz_9026;
  wire       [31:0]   _zz_9027;
  wire       [31:0]   _zz_9028;
  wire       [15:0]   _zz_9029;
  wire       [31:0]   _zz_9030;
  wire       [31:0]   _zz_9031;
  wire       [15:0]   _zz_9032;
  wire       [15:0]   _zz_9033;
  wire       [15:0]   _zz_9034;
  wire       [15:0]   _zz_9035;
  wire       [15:0]   _zz_9036;
  wire       [15:0]   _zz_9037;
  wire       [15:0]   _zz_9038;
  wire       [15:0]   _zz_9039;
  wire       [15:0]   _zz_9040;
  wire       [15:0]   _zz_9041;
  wire       [15:0]   _zz_9042;
  wire       [15:0]   _zz_9043;
  wire       [15:0]   _zz_9044;
  wire       [15:0]   _zz_9045;
  wire       [15:0]   _zz_9046;
  wire       [15:0]   _zz_9047;
  wire       [15:0]   _zz_9048;
  wire       [31:0]   _zz_9049;
  wire       [31:0]   _zz_9050;
  wire       [15:0]   _zz_9051;
  wire       [31:0]   _zz_9052;
  wire       [31:0]   _zz_9053;
  wire       [15:0]   _zz_9054;
  wire       [15:0]   _zz_9055;
  wire       [15:0]   _zz_9056;
  wire       [15:0]   _zz_9057;
  wire       [15:0]   _zz_9058;
  wire       [15:0]   _zz_9059;
  wire       [15:0]   _zz_9060;
  wire       [15:0]   _zz_9061;
  wire       [15:0]   _zz_9062;
  wire       [15:0]   _zz_9063;
  wire       [15:0]   _zz_9064;
  wire       [15:0]   _zz_9065;
  wire       [15:0]   _zz_9066;
  wire       [15:0]   _zz_9067;
  wire       [15:0]   _zz_9068;
  wire       [15:0]   _zz_9069;
  wire       [15:0]   _zz_9070;
  wire       [31:0]   _zz_9071;
  wire       [31:0]   _zz_9072;
  wire       [15:0]   _zz_9073;
  wire       [31:0]   _zz_9074;
  wire       [31:0]   _zz_9075;
  wire       [15:0]   _zz_9076;
  wire       [15:0]   _zz_9077;
  wire       [15:0]   _zz_9078;
  wire       [15:0]   _zz_9079;
  wire       [15:0]   _zz_9080;
  wire       [15:0]   _zz_9081;
  wire       [15:0]   _zz_9082;
  wire       [15:0]   _zz_9083;
  wire       [15:0]   _zz_9084;
  wire       [15:0]   _zz_9085;
  wire       [15:0]   _zz_9086;
  wire       [15:0]   _zz_9087;
  wire       [15:0]   _zz_9088;
  wire       [15:0]   _zz_9089;
  wire       [15:0]   _zz_9090;
  wire       [15:0]   _zz_9091;
  wire       [15:0]   _zz_9092;
  wire       [31:0]   _zz_9093;
  wire       [31:0]   _zz_9094;
  wire       [15:0]   _zz_9095;
  wire       [31:0]   _zz_9096;
  wire       [31:0]   _zz_9097;
  wire       [15:0]   _zz_9098;
  wire       [15:0]   _zz_9099;
  wire       [15:0]   _zz_9100;
  wire       [15:0]   _zz_9101;
  wire       [15:0]   _zz_9102;
  wire       [15:0]   _zz_9103;
  wire       [15:0]   _zz_9104;
  wire       [15:0]   _zz_9105;
  wire       [15:0]   _zz_9106;
  wire       [15:0]   _zz_9107;
  wire       [15:0]   _zz_9108;
  wire       [15:0]   _zz_9109;
  wire       [15:0]   _zz_9110;
  wire       [15:0]   _zz_9111;
  wire       [15:0]   _zz_9112;
  wire       [15:0]   _zz_9113;
  wire       [15:0]   _zz_9114;
  wire       [31:0]   _zz_9115;
  wire       [31:0]   _zz_9116;
  wire       [15:0]   _zz_9117;
  wire       [31:0]   _zz_9118;
  wire       [31:0]   _zz_9119;
  wire       [15:0]   _zz_9120;
  wire       [15:0]   _zz_9121;
  wire       [15:0]   _zz_9122;
  wire       [15:0]   _zz_9123;
  wire       [15:0]   _zz_9124;
  wire       [15:0]   _zz_9125;
  wire       [15:0]   _zz_9126;
  wire       [15:0]   _zz_9127;
  wire       [15:0]   _zz_9128;
  wire       [15:0]   _zz_9129;
  wire       [15:0]   _zz_9130;
  wire       [15:0]   _zz_9131;
  wire       [15:0]   _zz_9132;
  wire       [15:0]   _zz_9133;
  wire       [15:0]   _zz_9134;
  wire       [15:0]   _zz_9135;
  wire       [15:0]   _zz_9136;
  wire       [31:0]   _zz_9137;
  wire       [31:0]   _zz_9138;
  wire       [15:0]   _zz_9139;
  wire       [31:0]   _zz_9140;
  wire       [31:0]   _zz_9141;
  wire       [15:0]   _zz_9142;
  wire       [15:0]   _zz_9143;
  wire       [15:0]   _zz_9144;
  wire       [15:0]   _zz_9145;
  wire       [15:0]   _zz_9146;
  wire       [15:0]   _zz_9147;
  wire       [15:0]   _zz_9148;
  wire       [15:0]   _zz_9149;
  wire       [15:0]   _zz_9150;
  wire       [15:0]   _zz_9151;
  wire       [15:0]   _zz_9152;
  wire       [15:0]   _zz_9153;
  wire       [15:0]   _zz_9154;
  wire       [15:0]   _zz_9155;
  wire       [15:0]   _zz_9156;
  wire       [15:0]   _zz_9157;
  wire       [15:0]   _zz_9158;
  wire       [31:0]   _zz_9159;
  wire       [31:0]   _zz_9160;
  wire       [15:0]   _zz_9161;
  wire       [31:0]   _zz_9162;
  wire       [31:0]   _zz_9163;
  wire       [15:0]   _zz_9164;
  wire       [15:0]   _zz_9165;
  wire       [15:0]   _zz_9166;
  wire       [15:0]   _zz_9167;
  wire       [15:0]   _zz_9168;
  wire       [15:0]   _zz_9169;
  wire       [15:0]   _zz_9170;
  wire       [15:0]   _zz_9171;
  wire       [15:0]   _zz_9172;
  wire       [15:0]   _zz_9173;
  wire       [15:0]   _zz_9174;
  wire       [15:0]   _zz_9175;
  wire       [15:0]   _zz_9176;
  wire       [15:0]   _zz_9177;
  wire       [15:0]   _zz_9178;
  wire       [15:0]   _zz_9179;
  wire       [15:0]   _zz_9180;
  wire       [31:0]   _zz_9181;
  wire       [31:0]   _zz_9182;
  wire       [15:0]   _zz_9183;
  wire       [31:0]   _zz_9184;
  wire       [31:0]   _zz_9185;
  wire       [15:0]   _zz_9186;
  wire       [15:0]   _zz_9187;
  wire       [15:0]   _zz_9188;
  wire       [15:0]   _zz_9189;
  wire       [15:0]   _zz_9190;
  wire       [15:0]   _zz_9191;
  wire       [15:0]   _zz_9192;
  wire       [15:0]   _zz_9193;
  wire       [15:0]   _zz_9194;
  wire       [15:0]   _zz_9195;
  wire       [15:0]   _zz_9196;
  wire       [15:0]   _zz_9197;
  wire       [15:0]   _zz_9198;
  wire       [15:0]   _zz_9199;
  wire       [15:0]   _zz_9200;
  wire       [15:0]   _zz_9201;
  wire       [15:0]   _zz_9202;
  wire       [31:0]   _zz_9203;
  wire       [31:0]   _zz_9204;
  wire       [15:0]   _zz_9205;
  wire       [31:0]   _zz_9206;
  wire       [31:0]   _zz_9207;
  wire       [15:0]   _zz_9208;
  wire       [15:0]   _zz_9209;
  wire       [15:0]   _zz_9210;
  wire       [15:0]   _zz_9211;
  wire       [15:0]   _zz_9212;
  wire       [15:0]   _zz_9213;
  wire       [15:0]   _zz_9214;
  wire       [15:0]   _zz_9215;
  wire       [15:0]   _zz_9216;
  wire       [15:0]   _zz_9217;
  wire       [15:0]   _zz_9218;
  wire       [15:0]   _zz_9219;
  wire       [15:0]   _zz_9220;
  wire       [15:0]   _zz_9221;
  wire       [15:0]   _zz_9222;
  wire       [15:0]   _zz_9223;
  wire       [15:0]   _zz_9224;
  wire       [31:0]   _zz_9225;
  wire       [31:0]   _zz_9226;
  wire       [15:0]   _zz_9227;
  wire       [31:0]   _zz_9228;
  wire       [31:0]   _zz_9229;
  wire       [15:0]   _zz_9230;
  wire       [15:0]   _zz_9231;
  wire       [15:0]   _zz_9232;
  wire       [15:0]   _zz_9233;
  wire       [15:0]   _zz_9234;
  wire       [15:0]   _zz_9235;
  wire       [15:0]   _zz_9236;
  wire       [15:0]   _zz_9237;
  wire       [15:0]   _zz_9238;
  wire       [15:0]   _zz_9239;
  wire       [15:0]   _zz_9240;
  wire       [15:0]   _zz_9241;
  wire       [15:0]   _zz_9242;
  wire       [15:0]   _zz_9243;
  wire       [15:0]   _zz_9244;
  wire       [15:0]   _zz_9245;
  wire       [15:0]   _zz_9246;
  wire       [31:0]   _zz_9247;
  wire       [31:0]   _zz_9248;
  wire       [15:0]   _zz_9249;
  wire       [31:0]   _zz_9250;
  wire       [31:0]   _zz_9251;
  wire       [15:0]   _zz_9252;
  wire       [15:0]   _zz_9253;
  wire       [15:0]   _zz_9254;
  wire       [15:0]   _zz_9255;
  wire       [15:0]   _zz_9256;
  wire       [15:0]   _zz_9257;
  wire       [15:0]   _zz_9258;
  wire       [15:0]   _zz_9259;
  wire       [15:0]   _zz_9260;
  wire       [15:0]   _zz_9261;
  wire       [15:0]   _zz_9262;
  wire       [15:0]   _zz_9263;
  wire       [15:0]   _zz_9264;
  wire       [15:0]   _zz_9265;
  wire       [15:0]   _zz_9266;
  wire       [15:0]   _zz_9267;
  wire       [15:0]   _zz_9268;
  wire       [31:0]   _zz_9269;
  wire       [31:0]   _zz_9270;
  wire       [15:0]   _zz_9271;
  wire       [31:0]   _zz_9272;
  wire       [31:0]   _zz_9273;
  wire       [15:0]   _zz_9274;
  wire       [15:0]   _zz_9275;
  wire       [15:0]   _zz_9276;
  wire       [15:0]   _zz_9277;
  wire       [15:0]   _zz_9278;
  wire       [15:0]   _zz_9279;
  wire       [15:0]   _zz_9280;
  wire       [15:0]   _zz_9281;
  wire       [15:0]   _zz_9282;
  wire       [15:0]   _zz_9283;
  wire       [15:0]   _zz_9284;
  wire       [15:0]   _zz_9285;
  wire       [15:0]   _zz_9286;
  wire       [15:0]   _zz_9287;
  wire       [15:0]   _zz_9288;
  wire       [15:0]   _zz_9289;
  wire       [15:0]   _zz_9290;
  wire       [31:0]   _zz_9291;
  wire       [31:0]   _zz_9292;
  wire       [15:0]   _zz_9293;
  wire       [31:0]   _zz_9294;
  wire       [31:0]   _zz_9295;
  wire       [15:0]   _zz_9296;
  wire       [15:0]   _zz_9297;
  wire       [15:0]   _zz_9298;
  wire       [15:0]   _zz_9299;
  wire       [15:0]   _zz_9300;
  wire       [15:0]   _zz_9301;
  wire       [15:0]   _zz_9302;
  wire       [15:0]   _zz_9303;
  wire       [15:0]   _zz_9304;
  wire       [15:0]   _zz_9305;
  wire       [15:0]   _zz_9306;
  wire       [15:0]   _zz_9307;
  wire       [15:0]   _zz_9308;
  wire       [15:0]   _zz_9309;
  wire       [15:0]   _zz_9310;
  wire       [15:0]   _zz_9311;
  wire       [15:0]   _zz_9312;
  wire       [31:0]   _zz_9313;
  wire       [31:0]   _zz_9314;
  wire       [15:0]   _zz_9315;
  wire       [31:0]   _zz_9316;
  wire       [31:0]   _zz_9317;
  wire       [15:0]   _zz_9318;
  wire       [15:0]   _zz_9319;
  wire       [15:0]   _zz_9320;
  wire       [15:0]   _zz_9321;
  wire       [15:0]   _zz_9322;
  wire       [15:0]   _zz_9323;
  wire       [15:0]   _zz_9324;
  wire       [15:0]   _zz_9325;
  wire       [15:0]   _zz_9326;
  wire       [15:0]   _zz_9327;
  wire       [15:0]   _zz_9328;
  wire       [15:0]   _zz_9329;
  wire       [15:0]   _zz_9330;
  wire       [15:0]   _zz_9331;
  wire       [15:0]   _zz_9332;
  wire       [15:0]   _zz_9333;
  wire       [15:0]   _zz_9334;
  wire       [31:0]   _zz_9335;
  wire       [31:0]   _zz_9336;
  wire       [15:0]   _zz_9337;
  wire       [31:0]   _zz_9338;
  wire       [31:0]   _zz_9339;
  wire       [15:0]   _zz_9340;
  wire       [15:0]   _zz_9341;
  wire       [15:0]   _zz_9342;
  wire       [15:0]   _zz_9343;
  wire       [15:0]   _zz_9344;
  wire       [15:0]   _zz_9345;
  wire       [15:0]   _zz_9346;
  wire       [15:0]   _zz_9347;
  wire       [15:0]   _zz_9348;
  wire       [15:0]   _zz_9349;
  wire       [15:0]   _zz_9350;
  wire       [15:0]   _zz_9351;
  wire       [15:0]   _zz_9352;
  wire       [15:0]   _zz_9353;
  wire       [15:0]   _zz_9354;
  wire       [15:0]   _zz_9355;
  wire       [15:0]   _zz_9356;
  wire       [31:0]   _zz_9357;
  wire       [31:0]   _zz_9358;
  wire       [15:0]   _zz_9359;
  wire       [31:0]   _zz_9360;
  wire       [31:0]   _zz_9361;
  wire       [15:0]   _zz_9362;
  wire       [15:0]   _zz_9363;
  wire       [15:0]   _zz_9364;
  wire       [15:0]   _zz_9365;
  wire       [15:0]   _zz_9366;
  wire       [15:0]   _zz_9367;
  wire       [15:0]   _zz_9368;
  wire       [15:0]   _zz_9369;
  wire       [15:0]   _zz_9370;
  wire       [15:0]   _zz_9371;
  wire       [15:0]   _zz_9372;
  wire       [15:0]   _zz_9373;
  wire       [15:0]   _zz_9374;
  wire       [15:0]   _zz_9375;
  wire       [15:0]   _zz_9376;
  wire       [15:0]   _zz_9377;
  wire       [15:0]   _zz_9378;
  wire       [31:0]   _zz_9379;
  wire       [31:0]   _zz_9380;
  wire       [15:0]   _zz_9381;
  wire       [31:0]   _zz_9382;
  wire       [31:0]   _zz_9383;
  wire       [15:0]   _zz_9384;
  wire       [15:0]   _zz_9385;
  wire       [15:0]   _zz_9386;
  wire       [15:0]   _zz_9387;
  wire       [15:0]   _zz_9388;
  wire       [15:0]   _zz_9389;
  wire       [15:0]   _zz_9390;
  wire       [15:0]   _zz_9391;
  wire       [15:0]   _zz_9392;
  wire       [15:0]   _zz_9393;
  wire       [15:0]   _zz_9394;
  wire       [15:0]   _zz_9395;
  wire       [15:0]   _zz_9396;
  wire       [15:0]   _zz_9397;
  wire       [15:0]   _zz_9398;
  wire       [15:0]   _zz_9399;
  wire       [15:0]   _zz_9400;
  wire       [31:0]   _zz_9401;
  wire       [31:0]   _zz_9402;
  wire       [15:0]   _zz_9403;
  wire       [31:0]   _zz_9404;
  wire       [31:0]   _zz_9405;
  wire       [15:0]   _zz_9406;
  wire       [15:0]   _zz_9407;
  wire       [15:0]   _zz_9408;
  wire       [15:0]   _zz_9409;
  wire       [15:0]   _zz_9410;
  wire       [15:0]   _zz_9411;
  wire       [15:0]   _zz_9412;
  wire       [15:0]   _zz_9413;
  wire       [15:0]   _zz_9414;
  wire       [15:0]   _zz_9415;
  wire       [15:0]   _zz_9416;
  wire       [15:0]   _zz_9417;
  wire       [15:0]   _zz_9418;
  wire       [15:0]   _zz_9419;
  wire       [15:0]   _zz_9420;
  wire       [15:0]   _zz_9421;
  wire       [15:0]   _zz_9422;
  wire       [31:0]   _zz_9423;
  wire       [31:0]   _zz_9424;
  wire       [15:0]   _zz_9425;
  wire       [31:0]   _zz_9426;
  wire       [31:0]   _zz_9427;
  wire       [15:0]   _zz_9428;
  wire       [15:0]   _zz_9429;
  wire       [15:0]   _zz_9430;
  wire       [15:0]   _zz_9431;
  wire       [15:0]   _zz_9432;
  wire       [15:0]   _zz_9433;
  wire       [15:0]   _zz_9434;
  wire       [15:0]   _zz_9435;
  wire       [15:0]   _zz_9436;
  wire       [15:0]   _zz_9437;
  wire       [15:0]   _zz_9438;
  wire       [15:0]   _zz_9439;
  wire       [15:0]   _zz_9440;
  wire       [15:0]   _zz_9441;
  wire       [15:0]   _zz_9442;
  wire       [15:0]   _zz_9443;
  wire       [15:0]   _zz_9444;
  wire       [31:0]   _zz_9445;
  wire       [31:0]   _zz_9446;
  wire       [15:0]   _zz_9447;
  wire       [31:0]   _zz_9448;
  wire       [31:0]   _zz_9449;
  wire       [15:0]   _zz_9450;
  wire       [15:0]   _zz_9451;
  wire       [15:0]   _zz_9452;
  wire       [15:0]   _zz_9453;
  wire       [15:0]   _zz_9454;
  wire       [15:0]   _zz_9455;
  wire       [15:0]   _zz_9456;
  wire       [15:0]   _zz_9457;
  wire       [15:0]   _zz_9458;
  wire       [15:0]   _zz_9459;
  wire       [15:0]   _zz_9460;
  wire       [15:0]   _zz_9461;
  wire       [15:0]   _zz_9462;
  wire       [15:0]   _zz_9463;
  wire       [15:0]   _zz_9464;
  wire       [15:0]   _zz_9465;
  wire       [15:0]   _zz_9466;
  wire       [31:0]   _zz_9467;
  wire       [31:0]   _zz_9468;
  wire       [15:0]   _zz_9469;
  wire       [31:0]   _zz_9470;
  wire       [31:0]   _zz_9471;
  wire       [15:0]   _zz_9472;
  wire       [15:0]   _zz_9473;
  wire       [15:0]   _zz_9474;
  wire       [15:0]   _zz_9475;
  wire       [15:0]   _zz_9476;
  wire       [15:0]   _zz_9477;
  wire       [15:0]   _zz_9478;
  wire       [15:0]   _zz_9479;
  wire       [15:0]   _zz_9480;
  wire       [15:0]   _zz_9481;
  wire       [15:0]   _zz_9482;
  wire       [15:0]   _zz_9483;
  wire       [15:0]   _zz_9484;
  wire       [15:0]   _zz_9485;
  wire       [15:0]   _zz_9486;
  wire       [15:0]   _zz_9487;
  wire       [15:0]   _zz_9488;
  wire       [31:0]   _zz_9489;
  wire       [31:0]   _zz_9490;
  wire       [15:0]   _zz_9491;
  wire       [31:0]   _zz_9492;
  wire       [31:0]   _zz_9493;
  wire       [15:0]   _zz_9494;
  wire       [15:0]   _zz_9495;
  wire       [15:0]   _zz_9496;
  wire       [15:0]   _zz_9497;
  wire       [15:0]   _zz_9498;
  wire       [15:0]   _zz_9499;
  wire       [15:0]   _zz_9500;
  wire       [15:0]   _zz_9501;
  wire       [15:0]   _zz_9502;
  wire       [15:0]   _zz_9503;
  wire       [15:0]   _zz_9504;
  wire       [15:0]   _zz_9505;
  wire       [15:0]   _zz_9506;
  wire       [15:0]   _zz_9507;
  wire       [15:0]   _zz_9508;
  wire       [15:0]   _zz_9509;
  wire       [15:0]   _zz_9510;
  wire       [31:0]   _zz_9511;
  wire       [31:0]   _zz_9512;
  wire       [15:0]   _zz_9513;
  wire       [31:0]   _zz_9514;
  wire       [31:0]   _zz_9515;
  wire       [15:0]   _zz_9516;
  wire       [15:0]   _zz_9517;
  wire       [15:0]   _zz_9518;
  wire       [15:0]   _zz_9519;
  wire       [15:0]   _zz_9520;
  wire       [15:0]   _zz_9521;
  wire       [15:0]   _zz_9522;
  wire       [15:0]   _zz_9523;
  wire       [15:0]   _zz_9524;
  wire       [15:0]   _zz_9525;
  wire       [15:0]   _zz_9526;
  wire       [15:0]   _zz_9527;
  wire       [15:0]   _zz_9528;
  wire       [15:0]   _zz_9529;
  wire       [15:0]   _zz_9530;
  wire       [15:0]   _zz_9531;
  wire       [15:0]   _zz_9532;
  wire       [31:0]   _zz_9533;
  wire       [31:0]   _zz_9534;
  wire       [15:0]   _zz_9535;
  wire       [31:0]   _zz_9536;
  wire       [31:0]   _zz_9537;
  wire       [15:0]   _zz_9538;
  wire       [15:0]   _zz_9539;
  wire       [15:0]   _zz_9540;
  wire       [15:0]   _zz_9541;
  wire       [15:0]   _zz_9542;
  wire       [15:0]   _zz_9543;
  wire       [15:0]   _zz_9544;
  wire       [15:0]   _zz_9545;
  wire       [15:0]   _zz_9546;
  wire       [15:0]   _zz_9547;
  wire       [15:0]   _zz_9548;
  wire       [15:0]   _zz_9549;
  wire       [15:0]   _zz_9550;
  wire       [15:0]   _zz_9551;
  wire       [15:0]   _zz_9552;
  wire       [15:0]   _zz_9553;
  wire       [15:0]   _zz_9554;
  wire       [31:0]   _zz_9555;
  wire       [31:0]   _zz_9556;
  wire       [15:0]   _zz_9557;
  wire       [31:0]   _zz_9558;
  wire       [31:0]   _zz_9559;
  wire       [15:0]   _zz_9560;
  wire       [15:0]   _zz_9561;
  wire       [15:0]   _zz_9562;
  wire       [15:0]   _zz_9563;
  wire       [15:0]   _zz_9564;
  wire       [15:0]   _zz_9565;
  wire       [15:0]   _zz_9566;
  wire       [15:0]   _zz_9567;
  wire       [15:0]   _zz_9568;
  wire       [15:0]   _zz_9569;
  wire       [15:0]   _zz_9570;
  wire       [15:0]   _zz_9571;
  wire       [15:0]   _zz_9572;
  wire       [15:0]   _zz_9573;
  wire       [15:0]   _zz_9574;
  wire       [15:0]   _zz_9575;
  wire       [15:0]   _zz_9576;
  wire       [31:0]   _zz_9577;
  wire       [31:0]   _zz_9578;
  wire       [15:0]   _zz_9579;
  wire       [31:0]   _zz_9580;
  wire       [31:0]   _zz_9581;
  wire       [15:0]   _zz_9582;
  wire       [15:0]   _zz_9583;
  wire       [15:0]   _zz_9584;
  wire       [15:0]   _zz_9585;
  wire       [15:0]   _zz_9586;
  wire       [15:0]   _zz_9587;
  wire       [15:0]   _zz_9588;
  wire       [15:0]   _zz_9589;
  wire       [15:0]   _zz_9590;
  wire       [15:0]   _zz_9591;
  wire       [15:0]   _zz_9592;
  wire       [15:0]   _zz_9593;
  wire       [15:0]   _zz_9594;
  wire       [15:0]   _zz_9595;
  wire       [15:0]   _zz_9596;
  wire       [15:0]   _zz_9597;
  wire       [15:0]   _zz_9598;
  wire       [31:0]   _zz_9599;
  wire       [31:0]   _zz_9600;
  wire       [15:0]   _zz_9601;
  wire       [31:0]   _zz_9602;
  wire       [31:0]   _zz_9603;
  wire       [15:0]   _zz_9604;
  wire       [15:0]   _zz_9605;
  wire       [15:0]   _zz_9606;
  wire       [15:0]   _zz_9607;
  wire       [15:0]   _zz_9608;
  wire       [15:0]   _zz_9609;
  wire       [15:0]   _zz_9610;
  wire       [15:0]   _zz_9611;
  wire       [15:0]   _zz_9612;
  wire       [15:0]   _zz_9613;
  wire       [15:0]   _zz_9614;
  wire       [15:0]   _zz_9615;
  wire       [15:0]   _zz_9616;
  wire       [15:0]   _zz_9617;
  wire       [15:0]   _zz_9618;
  wire       [15:0]   _zz_9619;
  wire       [15:0]   _zz_9620;
  wire       [31:0]   _zz_9621;
  wire       [31:0]   _zz_9622;
  wire       [15:0]   _zz_9623;
  wire       [31:0]   _zz_9624;
  wire       [31:0]   _zz_9625;
  wire       [15:0]   _zz_9626;
  wire       [15:0]   _zz_9627;
  wire       [15:0]   _zz_9628;
  wire       [15:0]   _zz_9629;
  wire       [15:0]   _zz_9630;
  wire       [15:0]   _zz_9631;
  wire       [15:0]   _zz_9632;
  wire       [15:0]   _zz_9633;
  wire       [15:0]   _zz_9634;
  wire       [15:0]   _zz_9635;
  wire       [15:0]   _zz_9636;
  wire       [15:0]   _zz_9637;
  wire       [15:0]   _zz_9638;
  wire       [15:0]   _zz_9639;
  wire       [15:0]   _zz_9640;
  wire       [15:0]   _zz_9641;
  wire       [15:0]   _zz_9642;
  wire       [31:0]   _zz_9643;
  wire       [31:0]   _zz_9644;
  wire       [15:0]   _zz_9645;
  wire       [31:0]   _zz_9646;
  wire       [31:0]   _zz_9647;
  wire       [15:0]   _zz_9648;
  wire       [15:0]   _zz_9649;
  wire       [15:0]   _zz_9650;
  wire       [15:0]   _zz_9651;
  wire       [15:0]   _zz_9652;
  wire       [15:0]   _zz_9653;
  wire       [15:0]   _zz_9654;
  wire       [15:0]   _zz_9655;
  wire       [15:0]   _zz_9656;
  wire       [15:0]   _zz_9657;
  wire       [15:0]   _zz_9658;
  wire       [15:0]   _zz_9659;
  wire       [15:0]   _zz_9660;
  wire       [15:0]   _zz_9661;
  wire       [15:0]   _zz_9662;
  wire       [15:0]   _zz_9663;
  wire       [15:0]   _zz_9664;
  wire       [31:0]   _zz_9665;
  wire       [31:0]   _zz_9666;
  wire       [15:0]   _zz_9667;
  wire       [31:0]   _zz_9668;
  wire       [31:0]   _zz_9669;
  wire       [15:0]   _zz_9670;
  wire       [15:0]   _zz_9671;
  wire       [15:0]   _zz_9672;
  wire       [15:0]   _zz_9673;
  wire       [15:0]   _zz_9674;
  wire       [15:0]   _zz_9675;
  wire       [15:0]   _zz_9676;
  wire       [15:0]   _zz_9677;
  wire       [15:0]   _zz_9678;
  wire       [15:0]   _zz_9679;
  wire       [15:0]   _zz_9680;
  wire       [15:0]   _zz_9681;
  wire       [15:0]   _zz_9682;
  wire       [15:0]   _zz_9683;
  wire       [15:0]   _zz_9684;
  wire       [15:0]   _zz_9685;
  wire       [15:0]   _zz_9686;
  wire       [31:0]   _zz_9687;
  wire       [31:0]   _zz_9688;
  wire       [15:0]   _zz_9689;
  wire       [31:0]   _zz_9690;
  wire       [31:0]   _zz_9691;
  wire       [15:0]   _zz_9692;
  wire       [15:0]   _zz_9693;
  wire       [15:0]   _zz_9694;
  wire       [15:0]   _zz_9695;
  wire       [15:0]   _zz_9696;
  wire       [15:0]   _zz_9697;
  wire       [15:0]   _zz_9698;
  wire       [15:0]   _zz_9699;
  wire       [15:0]   _zz_9700;
  wire       [15:0]   _zz_9701;
  wire       [15:0]   _zz_9702;
  wire       [15:0]   _zz_9703;
  wire       [15:0]   _zz_9704;
  wire       [15:0]   _zz_9705;
  wire       [15:0]   _zz_9706;
  wire       [15:0]   _zz_9707;
  wire       [15:0]   _zz_9708;
  wire       [31:0]   _zz_9709;
  wire       [31:0]   _zz_9710;
  wire       [15:0]   _zz_9711;
  wire       [31:0]   _zz_9712;
  wire       [31:0]   _zz_9713;
  wire       [15:0]   _zz_9714;
  wire       [15:0]   _zz_9715;
  wire       [15:0]   _zz_9716;
  wire       [15:0]   _zz_9717;
  wire       [15:0]   _zz_9718;
  wire       [15:0]   _zz_9719;
  wire       [15:0]   _zz_9720;
  wire       [15:0]   _zz_9721;
  wire       [15:0]   _zz_9722;
  wire       [15:0]   _zz_9723;
  wire       [15:0]   _zz_9724;
  wire       [15:0]   _zz_9725;
  wire       [15:0]   _zz_9726;
  wire       [15:0]   _zz_9727;
  wire       [15:0]   _zz_9728;
  wire       [15:0]   _zz_9729;
  wire       [15:0]   _zz_9730;
  wire       [31:0]   _zz_9731;
  wire       [31:0]   _zz_9732;
  wire       [15:0]   _zz_9733;
  wire       [31:0]   _zz_9734;
  wire       [31:0]   _zz_9735;
  wire       [15:0]   _zz_9736;
  wire       [15:0]   _zz_9737;
  wire       [15:0]   _zz_9738;
  wire       [15:0]   _zz_9739;
  wire       [15:0]   _zz_9740;
  wire       [15:0]   _zz_9741;
  wire       [15:0]   _zz_9742;
  wire       [15:0]   _zz_9743;
  wire       [15:0]   _zz_9744;
  wire       [15:0]   _zz_9745;
  wire       [15:0]   _zz_9746;
  wire       [15:0]   _zz_9747;
  wire       [15:0]   _zz_9748;
  wire       [15:0]   _zz_9749;
  wire       [15:0]   _zz_9750;
  wire       [15:0]   _zz_9751;
  wire       [15:0]   _zz_9752;
  wire       [31:0]   _zz_9753;
  wire       [31:0]   _zz_9754;
  wire       [15:0]   _zz_9755;
  wire       [31:0]   _zz_9756;
  wire       [31:0]   _zz_9757;
  wire       [15:0]   _zz_9758;
  wire       [15:0]   _zz_9759;
  wire       [15:0]   _zz_9760;
  wire       [15:0]   _zz_9761;
  wire       [15:0]   _zz_9762;
  wire       [15:0]   _zz_9763;
  wire       [15:0]   _zz_9764;
  wire       [15:0]   _zz_9765;
  wire       [15:0]   _zz_9766;
  wire       [15:0]   _zz_9767;
  wire       [15:0]   _zz_9768;
  wire       [15:0]   _zz_9769;
  wire       [15:0]   _zz_9770;
  wire       [15:0]   _zz_9771;
  wire       [15:0]   _zz_9772;
  wire       [15:0]   _zz_9773;
  wire       [15:0]   _zz_9774;
  wire       [31:0]   _zz_9775;
  wire       [31:0]   _zz_9776;
  wire       [15:0]   _zz_9777;
  wire       [31:0]   _zz_9778;
  wire       [31:0]   _zz_9779;
  wire       [15:0]   _zz_9780;
  wire       [15:0]   _zz_9781;
  wire       [15:0]   _zz_9782;
  wire       [15:0]   _zz_9783;
  wire       [15:0]   _zz_9784;
  wire       [15:0]   _zz_9785;
  wire       [15:0]   _zz_9786;
  wire       [15:0]   _zz_9787;
  wire       [15:0]   _zz_9788;
  wire       [15:0]   _zz_9789;
  wire       [15:0]   _zz_9790;
  wire       [15:0]   _zz_9791;
  wire       [15:0]   _zz_9792;
  wire       [15:0]   _zz_9793;
  wire       [15:0]   _zz_9794;
  wire       [15:0]   _zz_9795;
  wire       [15:0]   _zz_9796;
  wire       [31:0]   _zz_9797;
  wire       [31:0]   _zz_9798;
  wire       [15:0]   _zz_9799;
  wire       [31:0]   _zz_9800;
  wire       [31:0]   _zz_9801;
  wire       [15:0]   _zz_9802;
  wire       [15:0]   _zz_9803;
  wire       [15:0]   _zz_9804;
  wire       [15:0]   _zz_9805;
  wire       [15:0]   _zz_9806;
  wire       [15:0]   _zz_9807;
  wire       [15:0]   _zz_9808;
  wire       [15:0]   _zz_9809;
  wire       [15:0]   _zz_9810;
  wire       [15:0]   _zz_9811;
  wire       [15:0]   _zz_9812;
  wire       [15:0]   _zz_9813;
  wire       [15:0]   _zz_9814;
  wire       [15:0]   _zz_9815;
  wire       [15:0]   _zz_9816;
  wire       [15:0]   _zz_9817;
  wire       [15:0]   _zz_9818;
  wire       [31:0]   _zz_9819;
  wire       [31:0]   _zz_9820;
  wire       [15:0]   _zz_9821;
  wire       [31:0]   _zz_9822;
  wire       [31:0]   _zz_9823;
  wire       [15:0]   _zz_9824;
  wire       [15:0]   _zz_9825;
  wire       [15:0]   _zz_9826;
  wire       [15:0]   _zz_9827;
  wire       [15:0]   _zz_9828;
  wire       [15:0]   _zz_9829;
  wire       [15:0]   _zz_9830;
  wire       [15:0]   _zz_9831;
  wire       [15:0]   _zz_9832;
  wire       [15:0]   _zz_9833;
  wire       [15:0]   _zz_9834;
  wire       [15:0]   _zz_9835;
  wire       [15:0]   _zz_9836;
  wire       [15:0]   _zz_9837;
  wire       [15:0]   _zz_9838;
  wire       [15:0]   _zz_9839;
  wire       [15:0]   _zz_9840;
  wire       [31:0]   _zz_9841;
  wire       [31:0]   _zz_9842;
  wire       [15:0]   _zz_9843;
  wire       [31:0]   _zz_9844;
  wire       [31:0]   _zz_9845;
  wire       [15:0]   _zz_9846;
  wire       [15:0]   _zz_9847;
  wire       [15:0]   _zz_9848;
  wire       [15:0]   _zz_9849;
  wire       [15:0]   _zz_9850;
  wire       [15:0]   _zz_9851;
  wire       [15:0]   _zz_9852;
  wire       [15:0]   _zz_9853;
  wire       [15:0]   _zz_9854;
  wire       [15:0]   _zz_9855;
  wire       [15:0]   _zz_9856;
  wire       [15:0]   _zz_9857;
  wire       [15:0]   _zz_9858;
  wire       [15:0]   _zz_9859;
  wire       [15:0]   _zz_9860;
  wire       [15:0]   _zz_9861;
  wire       [15:0]   _zz_9862;
  wire       [31:0]   _zz_9863;
  wire       [31:0]   _zz_9864;
  wire       [15:0]   _zz_9865;
  wire       [31:0]   _zz_9866;
  wire       [31:0]   _zz_9867;
  wire       [15:0]   _zz_9868;
  wire       [15:0]   _zz_9869;
  wire       [15:0]   _zz_9870;
  wire       [15:0]   _zz_9871;
  wire       [15:0]   _zz_9872;
  wire       [15:0]   _zz_9873;
  wire       [15:0]   _zz_9874;
  wire       [15:0]   _zz_9875;
  wire       [15:0]   _zz_9876;
  wire       [15:0]   _zz_9877;
  wire       [15:0]   _zz_9878;
  wire       [15:0]   _zz_9879;
  wire       [15:0]   _zz_9880;
  wire       [15:0]   _zz_9881;
  wire       [15:0]   _zz_9882;
  wire       [15:0]   _zz_9883;
  wire       [15:0]   _zz_9884;
  wire       [31:0]   _zz_9885;
  wire       [31:0]   _zz_9886;
  wire       [15:0]   _zz_9887;
  wire       [31:0]   _zz_9888;
  wire       [31:0]   _zz_9889;
  wire       [15:0]   _zz_9890;
  wire       [15:0]   _zz_9891;
  wire       [15:0]   _zz_9892;
  wire       [15:0]   _zz_9893;
  wire       [15:0]   _zz_9894;
  wire       [15:0]   _zz_9895;
  wire       [15:0]   _zz_9896;
  wire       [15:0]   _zz_9897;
  wire       [15:0]   _zz_9898;
  wire       [15:0]   _zz_9899;
  wire       [15:0]   _zz_9900;
  wire       [15:0]   _zz_9901;
  wire       [15:0]   _zz_9902;
  wire       [15:0]   _zz_9903;
  wire       [15:0]   _zz_9904;
  wire       [15:0]   _zz_9905;
  wire       [15:0]   _zz_9906;
  wire       [31:0]   _zz_9907;
  wire       [31:0]   _zz_9908;
  wire       [15:0]   _zz_9909;
  wire       [31:0]   _zz_9910;
  wire       [31:0]   _zz_9911;
  wire       [15:0]   _zz_9912;
  wire       [15:0]   _zz_9913;
  wire       [15:0]   _zz_9914;
  wire       [15:0]   _zz_9915;
  wire       [15:0]   _zz_9916;
  wire       [15:0]   _zz_9917;
  wire       [15:0]   _zz_9918;
  wire       [15:0]   _zz_9919;
  wire       [15:0]   _zz_9920;
  wire       [15:0]   _zz_9921;
  wire       [15:0]   _zz_9922;
  wire       [15:0]   _zz_9923;
  wire       [15:0]   _zz_9924;
  wire       [15:0]   _zz_9925;
  wire       [15:0]   _zz_9926;
  wire       [15:0]   _zz_9927;
  wire       [15:0]   _zz_9928;
  wire       [31:0]   _zz_9929;
  wire       [31:0]   _zz_9930;
  wire       [15:0]   _zz_9931;
  wire       [31:0]   _zz_9932;
  wire       [31:0]   _zz_9933;
  wire       [15:0]   _zz_9934;
  wire       [15:0]   _zz_9935;
  wire       [15:0]   _zz_9936;
  wire       [15:0]   _zz_9937;
  wire       [15:0]   _zz_9938;
  wire       [15:0]   _zz_9939;
  wire       [15:0]   _zz_9940;
  wire       [15:0]   _zz_9941;
  wire       [15:0]   _zz_9942;
  wire       [15:0]   _zz_9943;
  wire       [15:0]   _zz_9944;
  wire       [15:0]   _zz_9945;
  wire       [15:0]   _zz_9946;
  wire       [15:0]   _zz_9947;
  wire       [15:0]   _zz_9948;
  wire       [15:0]   _zz_9949;
  wire       [15:0]   _zz_9950;
  wire       [31:0]   _zz_9951;
  wire       [31:0]   _zz_9952;
  wire       [15:0]   _zz_9953;
  wire       [31:0]   _zz_9954;
  wire       [31:0]   _zz_9955;
  wire       [15:0]   _zz_9956;
  wire       [15:0]   _zz_9957;
  wire       [15:0]   _zz_9958;
  wire       [15:0]   _zz_9959;
  wire       [15:0]   _zz_9960;
  wire       [15:0]   _zz_9961;
  wire       [15:0]   _zz_9962;
  wire       [15:0]   _zz_9963;
  wire       [15:0]   _zz_9964;
  wire       [15:0]   _zz_9965;
  wire       [15:0]   _zz_9966;
  wire       [15:0]   _zz_9967;
  wire       [15:0]   _zz_9968;
  wire       [15:0]   _zz_9969;
  wire       [15:0]   _zz_9970;
  wire       [15:0]   _zz_9971;
  wire       [15:0]   _zz_9972;
  wire       [31:0]   _zz_9973;
  wire       [31:0]   _zz_9974;
  wire       [15:0]   _zz_9975;
  wire       [31:0]   _zz_9976;
  wire       [31:0]   _zz_9977;
  wire       [15:0]   _zz_9978;
  wire       [15:0]   _zz_9979;
  wire       [15:0]   _zz_9980;
  wire       [15:0]   _zz_9981;
  wire       [15:0]   _zz_9982;
  wire       [15:0]   _zz_9983;
  wire       [15:0]   _zz_9984;
  wire       [15:0]   _zz_9985;
  wire       [15:0]   _zz_9986;
  wire       [15:0]   _zz_9987;
  wire       [15:0]   _zz_9988;
  wire       [15:0]   _zz_9989;
  wire       [15:0]   _zz_9990;
  wire       [15:0]   _zz_9991;
  wire       [15:0]   _zz_9992;
  wire       [15:0]   _zz_9993;
  wire       [15:0]   _zz_9994;
  wire       [31:0]   _zz_9995;
  wire       [31:0]   _zz_9996;
  wire       [15:0]   _zz_9997;
  wire       [31:0]   _zz_9998;
  wire       [31:0]   _zz_9999;
  wire       [15:0]   _zz_10000;
  wire       [15:0]   _zz_10001;
  wire       [15:0]   _zz_10002;
  wire       [15:0]   _zz_10003;
  wire       [15:0]   _zz_10004;
  wire       [15:0]   _zz_10005;
  wire       [15:0]   _zz_10006;
  wire       [15:0]   _zz_10007;
  wire       [15:0]   _zz_10008;
  wire       [15:0]   _zz_10009;
  wire       [15:0]   _zz_10010;
  wire       [15:0]   _zz_10011;
  wire       [15:0]   _zz_10012;
  wire       [15:0]   _zz_10013;
  wire       [15:0]   _zz_10014;
  wire       [15:0]   _zz_10015;
  wire       [15:0]   _zz_10016;
  wire       [31:0]   _zz_10017;
  wire       [31:0]   _zz_10018;
  wire       [15:0]   _zz_10019;
  wire       [31:0]   _zz_10020;
  wire       [31:0]   _zz_10021;
  wire       [15:0]   _zz_10022;
  wire       [15:0]   _zz_10023;
  wire       [15:0]   _zz_10024;
  wire       [15:0]   _zz_10025;
  wire       [15:0]   _zz_10026;
  wire       [15:0]   _zz_10027;
  wire       [15:0]   _zz_10028;
  wire       [15:0]   _zz_10029;
  wire       [15:0]   _zz_10030;
  wire       [15:0]   _zz_10031;
  wire       [15:0]   _zz_10032;
  wire       [15:0]   _zz_10033;
  wire       [15:0]   _zz_10034;
  wire       [15:0]   _zz_10035;
  wire       [15:0]   _zz_10036;
  wire       [15:0]   _zz_10037;
  wire       [15:0]   _zz_10038;
  wire       [31:0]   _zz_10039;
  wire       [31:0]   _zz_10040;
  wire       [15:0]   _zz_10041;
  wire       [31:0]   _zz_10042;
  wire       [31:0]   _zz_10043;
  wire       [15:0]   _zz_10044;
  wire       [15:0]   _zz_10045;
  wire       [15:0]   _zz_10046;
  wire       [15:0]   _zz_10047;
  wire       [15:0]   _zz_10048;
  wire       [15:0]   _zz_10049;
  wire       [15:0]   _zz_10050;
  wire       [15:0]   _zz_10051;
  wire       [15:0]   _zz_10052;
  wire       [15:0]   _zz_10053;
  wire       [15:0]   _zz_10054;
  wire       [15:0]   _zz_10055;
  wire       [15:0]   _zz_10056;
  wire       [15:0]   _zz_10057;
  wire       [15:0]   _zz_10058;
  wire       [15:0]   _zz_10059;
  wire       [15:0]   _zz_10060;
  wire       [31:0]   _zz_10061;
  wire       [31:0]   _zz_10062;
  wire       [15:0]   _zz_10063;
  wire       [31:0]   _zz_10064;
  wire       [31:0]   _zz_10065;
  wire       [15:0]   _zz_10066;
  wire       [15:0]   _zz_10067;
  wire       [15:0]   _zz_10068;
  wire       [15:0]   _zz_10069;
  wire       [15:0]   _zz_10070;
  wire       [15:0]   _zz_10071;
  wire       [15:0]   _zz_10072;
  wire       [15:0]   _zz_10073;
  wire       [15:0]   _zz_10074;
  wire       [15:0]   _zz_10075;
  wire       [15:0]   _zz_10076;
  wire       [15:0]   _zz_10077;
  wire       [15:0]   _zz_10078;
  wire       [15:0]   _zz_10079;
  wire       [15:0]   _zz_10080;
  wire       [15:0]   _zz_10081;
  wire       [15:0]   _zz_10082;
  wire       [31:0]   _zz_10083;
  wire       [31:0]   _zz_10084;
  wire       [15:0]   _zz_10085;
  wire       [31:0]   _zz_10086;
  wire       [31:0]   _zz_10087;
  wire       [15:0]   _zz_10088;
  wire       [15:0]   _zz_10089;
  wire       [15:0]   _zz_10090;
  wire       [15:0]   _zz_10091;
  wire       [15:0]   _zz_10092;
  wire       [15:0]   _zz_10093;
  wire       [15:0]   _zz_10094;
  wire       [15:0]   _zz_10095;
  wire       [15:0]   _zz_10096;
  wire       [15:0]   _zz_10097;
  wire       [15:0]   _zz_10098;
  wire       [15:0]   _zz_10099;
  wire       [15:0]   _zz_10100;
  wire       [15:0]   _zz_10101;
  wire       [15:0]   _zz_10102;
  wire       [15:0]   _zz_10103;
  wire       [15:0]   _zz_10104;
  wire       [31:0]   _zz_10105;
  wire       [31:0]   _zz_10106;
  wire       [15:0]   _zz_10107;
  wire       [31:0]   _zz_10108;
  wire       [31:0]   _zz_10109;
  wire       [15:0]   _zz_10110;
  wire       [15:0]   _zz_10111;
  wire       [15:0]   _zz_10112;
  wire       [15:0]   _zz_10113;
  wire       [15:0]   _zz_10114;
  wire       [15:0]   _zz_10115;
  wire       [15:0]   _zz_10116;
  wire       [15:0]   _zz_10117;
  wire       [15:0]   _zz_10118;
  wire       [15:0]   _zz_10119;
  wire       [15:0]   _zz_10120;
  wire       [15:0]   _zz_10121;
  wire       [15:0]   _zz_10122;
  wire       [15:0]   _zz_10123;
  wire       [15:0]   _zz_10124;
  wire       [15:0]   _zz_10125;
  wire       [15:0]   _zz_10126;
  wire       [31:0]   _zz_10127;
  wire       [31:0]   _zz_10128;
  wire       [15:0]   _zz_10129;
  wire       [31:0]   _zz_10130;
  wire       [31:0]   _zz_10131;
  wire       [15:0]   _zz_10132;
  wire       [15:0]   _zz_10133;
  wire       [15:0]   _zz_10134;
  wire       [15:0]   _zz_10135;
  wire       [15:0]   _zz_10136;
  wire       [15:0]   _zz_10137;
  wire       [15:0]   _zz_10138;
  wire       [15:0]   _zz_10139;
  wire       [15:0]   _zz_10140;
  wire       [15:0]   _zz_10141;
  wire       [15:0]   _zz_10142;
  wire       [15:0]   _zz_10143;
  wire       [15:0]   _zz_10144;
  wire       [15:0]   _zz_10145;
  wire       [15:0]   _zz_10146;
  wire       [15:0]   _zz_10147;
  wire       [15:0]   _zz_10148;
  wire       [31:0]   _zz_10149;
  wire       [31:0]   _zz_10150;
  wire       [15:0]   _zz_10151;
  wire       [31:0]   _zz_10152;
  wire       [31:0]   _zz_10153;
  wire       [15:0]   _zz_10154;
  wire       [15:0]   _zz_10155;
  wire       [15:0]   _zz_10156;
  wire       [15:0]   _zz_10157;
  wire       [15:0]   _zz_10158;
  wire       [15:0]   _zz_10159;
  wire       [15:0]   _zz_10160;
  wire       [15:0]   _zz_10161;
  wire       [15:0]   _zz_10162;
  wire       [15:0]   _zz_10163;
  wire       [15:0]   _zz_10164;
  wire       [15:0]   _zz_10165;
  wire       [15:0]   _zz_10166;
  wire       [15:0]   _zz_10167;
  wire       [15:0]   _zz_10168;
  wire       [15:0]   _zz_10169;
  wire       [15:0]   _zz_10170;
  wire       [31:0]   _zz_10171;
  wire       [31:0]   _zz_10172;
  wire       [15:0]   _zz_10173;
  wire       [31:0]   _zz_10174;
  wire       [31:0]   _zz_10175;
  wire       [15:0]   _zz_10176;
  wire       [15:0]   _zz_10177;
  wire       [15:0]   _zz_10178;
  wire       [15:0]   _zz_10179;
  wire       [15:0]   _zz_10180;
  wire       [15:0]   _zz_10181;
  wire       [15:0]   _zz_10182;
  wire       [15:0]   _zz_10183;
  wire       [15:0]   _zz_10184;
  wire       [15:0]   _zz_10185;
  wire       [15:0]   _zz_10186;
  wire       [15:0]   _zz_10187;
  wire       [15:0]   _zz_10188;
  wire       [15:0]   _zz_10189;
  wire       [15:0]   _zz_10190;
  wire       [15:0]   _zz_10191;
  wire       [15:0]   _zz_10192;
  wire       [31:0]   _zz_10193;
  wire       [31:0]   _zz_10194;
  wire       [15:0]   _zz_10195;
  wire       [31:0]   _zz_10196;
  wire       [31:0]   _zz_10197;
  wire       [15:0]   _zz_10198;
  wire       [15:0]   _zz_10199;
  wire       [15:0]   _zz_10200;
  wire       [15:0]   _zz_10201;
  wire       [15:0]   _zz_10202;
  wire       [15:0]   _zz_10203;
  wire       [15:0]   _zz_10204;
  wire       [15:0]   _zz_10205;
  wire       [15:0]   _zz_10206;
  wire       [15:0]   _zz_10207;
  wire       [15:0]   _zz_10208;
  wire       [15:0]   _zz_10209;
  wire       [15:0]   _zz_10210;
  wire       [15:0]   _zz_10211;
  wire       [15:0]   _zz_10212;
  wire       [15:0]   _zz_10213;
  wire       [15:0]   _zz_10214;
  wire       [31:0]   _zz_10215;
  wire       [31:0]   _zz_10216;
  wire       [15:0]   _zz_10217;
  wire       [31:0]   _zz_10218;
  wire       [31:0]   _zz_10219;
  wire       [15:0]   _zz_10220;
  wire       [15:0]   _zz_10221;
  wire       [15:0]   _zz_10222;
  wire       [15:0]   _zz_10223;
  wire       [15:0]   _zz_10224;
  wire       [15:0]   _zz_10225;
  wire       [15:0]   _zz_10226;
  wire       [15:0]   _zz_10227;
  wire       [15:0]   _zz_10228;
  wire       [15:0]   _zz_10229;
  wire       [15:0]   _zz_10230;
  wire       [15:0]   _zz_10231;
  wire       [15:0]   _zz_10232;
  wire       [15:0]   _zz_10233;
  wire       [15:0]   _zz_10234;
  wire       [15:0]   _zz_10235;
  wire       [15:0]   _zz_10236;
  wire       [31:0]   _zz_10237;
  wire       [31:0]   _zz_10238;
  wire       [15:0]   _zz_10239;
  wire       [31:0]   _zz_10240;
  wire       [31:0]   _zz_10241;
  wire       [15:0]   _zz_10242;
  wire       [15:0]   _zz_10243;
  wire       [15:0]   _zz_10244;
  wire       [15:0]   _zz_10245;
  wire       [15:0]   _zz_10246;
  wire       [15:0]   _zz_10247;
  wire       [15:0]   _zz_10248;
  wire       [15:0]   _zz_10249;
  wire       [15:0]   _zz_10250;
  wire       [15:0]   _zz_10251;
  wire       [15:0]   _zz_10252;
  wire       [15:0]   _zz_10253;
  wire       [15:0]   _zz_10254;
  wire       [15:0]   _zz_10255;
  wire       [15:0]   _zz_10256;
  wire       [15:0]   _zz_10257;
  wire       [15:0]   _zz_10258;
  wire       [31:0]   _zz_10259;
  wire       [31:0]   _zz_10260;
  wire       [15:0]   _zz_10261;
  wire       [31:0]   _zz_10262;
  wire       [31:0]   _zz_10263;
  wire       [15:0]   _zz_10264;
  wire       [15:0]   _zz_10265;
  wire       [15:0]   _zz_10266;
  wire       [15:0]   _zz_10267;
  wire       [15:0]   _zz_10268;
  wire       [15:0]   _zz_10269;
  wire       [15:0]   _zz_10270;
  wire       [15:0]   _zz_10271;
  wire       [15:0]   _zz_10272;
  wire       [15:0]   _zz_10273;
  wire       [15:0]   _zz_10274;
  wire       [15:0]   _zz_10275;
  wire       [15:0]   _zz_10276;
  wire       [15:0]   _zz_10277;
  wire       [15:0]   _zz_10278;
  wire       [15:0]   _zz_10279;
  wire       [15:0]   _zz_10280;
  wire       [31:0]   _zz_10281;
  wire       [31:0]   _zz_10282;
  wire       [15:0]   _zz_10283;
  wire       [31:0]   _zz_10284;
  wire       [31:0]   _zz_10285;
  wire       [15:0]   _zz_10286;
  wire       [15:0]   _zz_10287;
  wire       [15:0]   _zz_10288;
  wire       [15:0]   _zz_10289;
  wire       [15:0]   _zz_10290;
  wire       [15:0]   _zz_10291;
  wire       [15:0]   _zz_10292;
  wire       [15:0]   _zz_10293;
  wire       [15:0]   _zz_10294;
  wire       [15:0]   _zz_10295;
  wire       [15:0]   _zz_10296;
  wire       [15:0]   _zz_10297;
  wire       [15:0]   _zz_10298;
  wire       [15:0]   _zz_10299;
  wire       [15:0]   _zz_10300;
  wire       [15:0]   _zz_10301;
  wire       [15:0]   _zz_10302;
  wire       [31:0]   _zz_10303;
  wire       [31:0]   _zz_10304;
  wire       [15:0]   _zz_10305;
  wire       [31:0]   _zz_10306;
  wire       [31:0]   _zz_10307;
  wire       [15:0]   _zz_10308;
  wire       [15:0]   _zz_10309;
  wire       [15:0]   _zz_10310;
  wire       [15:0]   _zz_10311;
  wire       [15:0]   _zz_10312;
  wire       [15:0]   _zz_10313;
  wire       [15:0]   _zz_10314;
  wire       [15:0]   _zz_10315;
  wire       [15:0]   _zz_10316;
  wire       [15:0]   _zz_10317;
  wire       [15:0]   _zz_10318;
  wire       [15:0]   _zz_10319;
  wire       [15:0]   _zz_10320;
  wire       [15:0]   _zz_10321;
  wire       [15:0]   _zz_10322;
  wire       [15:0]   _zz_10323;
  wire       [15:0]   _zz_10324;
  wire       [31:0]   _zz_10325;
  wire       [31:0]   _zz_10326;
  wire       [15:0]   _zz_10327;
  wire       [31:0]   _zz_10328;
  wire       [31:0]   _zz_10329;
  wire       [15:0]   _zz_10330;
  wire       [15:0]   _zz_10331;
  wire       [15:0]   _zz_10332;
  wire       [15:0]   _zz_10333;
  wire       [15:0]   _zz_10334;
  wire       [15:0]   _zz_10335;
  wire       [15:0]   _zz_10336;
  wire       [15:0]   _zz_10337;
  wire       [15:0]   _zz_10338;
  wire       [15:0]   _zz_10339;
  wire       [15:0]   _zz_10340;
  wire       [15:0]   _zz_10341;
  wire       [15:0]   _zz_10342;
  wire       [15:0]   _zz_10343;
  wire       [15:0]   _zz_10344;
  wire       [15:0]   _zz_10345;
  wire       [15:0]   _zz_10346;
  wire       [31:0]   _zz_10347;
  wire       [31:0]   _zz_10348;
  wire       [15:0]   _zz_10349;
  wire       [31:0]   _zz_10350;
  wire       [31:0]   _zz_10351;
  wire       [15:0]   _zz_10352;
  wire       [15:0]   _zz_10353;
  wire       [15:0]   _zz_10354;
  wire       [15:0]   _zz_10355;
  wire       [15:0]   _zz_10356;
  wire       [15:0]   _zz_10357;
  wire       [15:0]   _zz_10358;
  wire       [15:0]   _zz_10359;
  wire       [15:0]   _zz_10360;
  wire       [15:0]   _zz_10361;
  wire       [15:0]   _zz_10362;
  wire       [15:0]   _zz_10363;
  wire       [15:0]   _zz_10364;
  wire       [15:0]   _zz_10365;
  wire       [15:0]   _zz_10366;
  wire       [15:0]   _zz_10367;
  wire       [15:0]   _zz_10368;
  wire       [31:0]   _zz_10369;
  wire       [31:0]   _zz_10370;
  wire       [15:0]   _zz_10371;
  wire       [31:0]   _zz_10372;
  wire       [31:0]   _zz_10373;
  wire       [15:0]   _zz_10374;
  wire       [15:0]   _zz_10375;
  wire       [15:0]   _zz_10376;
  wire       [15:0]   _zz_10377;
  wire       [15:0]   _zz_10378;
  wire       [15:0]   _zz_10379;
  wire       [15:0]   _zz_10380;
  wire       [15:0]   _zz_10381;
  wire       [15:0]   _zz_10382;
  wire       [15:0]   _zz_10383;
  wire       [15:0]   _zz_10384;
  wire       [15:0]   _zz_10385;
  wire       [15:0]   _zz_10386;
  wire       [15:0]   _zz_10387;
  wire       [15:0]   _zz_10388;
  wire       [15:0]   _zz_10389;
  wire       [15:0]   _zz_10390;
  wire       [31:0]   _zz_10391;
  wire       [31:0]   _zz_10392;
  wire       [15:0]   _zz_10393;
  wire       [31:0]   _zz_10394;
  wire       [31:0]   _zz_10395;
  wire       [15:0]   _zz_10396;
  wire       [15:0]   _zz_10397;
  wire       [15:0]   _zz_10398;
  wire       [15:0]   _zz_10399;
  wire       [15:0]   _zz_10400;
  wire       [15:0]   _zz_10401;
  wire       [15:0]   _zz_10402;
  wire       [15:0]   _zz_10403;
  wire       [15:0]   _zz_10404;
  wire       [15:0]   _zz_10405;
  wire       [15:0]   _zz_10406;
  wire       [15:0]   _zz_10407;
  wire       [15:0]   _zz_10408;
  wire       [15:0]   _zz_10409;
  wire       [15:0]   _zz_10410;
  wire       [15:0]   _zz_10411;
  wire       [15:0]   _zz_10412;
  wire       [31:0]   _zz_10413;
  wire       [31:0]   _zz_10414;
  wire       [15:0]   _zz_10415;
  wire       [31:0]   _zz_10416;
  wire       [31:0]   _zz_10417;
  wire       [15:0]   _zz_10418;
  wire       [15:0]   _zz_10419;
  wire       [15:0]   _zz_10420;
  wire       [15:0]   _zz_10421;
  wire       [15:0]   _zz_10422;
  wire       [15:0]   _zz_10423;
  wire       [15:0]   _zz_10424;
  wire       [15:0]   _zz_10425;
  wire       [15:0]   _zz_10426;
  wire       [15:0]   _zz_10427;
  wire       [15:0]   _zz_10428;
  wire       [15:0]   _zz_10429;
  wire       [15:0]   _zz_10430;
  wire       [15:0]   _zz_10431;
  wire       [15:0]   _zz_10432;
  wire       [15:0]   _zz_10433;
  wire       [15:0]   _zz_10434;
  wire       [31:0]   _zz_10435;
  wire       [31:0]   _zz_10436;
  wire       [15:0]   _zz_10437;
  wire       [31:0]   _zz_10438;
  wire       [31:0]   _zz_10439;
  wire       [15:0]   _zz_10440;
  wire       [15:0]   _zz_10441;
  wire       [15:0]   _zz_10442;
  wire       [15:0]   _zz_10443;
  wire       [15:0]   _zz_10444;
  wire       [15:0]   _zz_10445;
  wire       [15:0]   _zz_10446;
  wire       [15:0]   _zz_10447;
  wire       [15:0]   _zz_10448;
  wire       [15:0]   _zz_10449;
  wire       [15:0]   _zz_10450;
  wire       [15:0]   _zz_10451;
  wire       [15:0]   _zz_10452;
  wire       [15:0]   _zz_10453;
  wire       [15:0]   _zz_10454;
  wire       [15:0]   _zz_10455;
  wire       [15:0]   _zz_10456;
  wire       [31:0]   _zz_10457;
  wire       [31:0]   _zz_10458;
  wire       [15:0]   _zz_10459;
  wire       [31:0]   _zz_10460;
  wire       [31:0]   _zz_10461;
  wire       [15:0]   _zz_10462;
  wire       [15:0]   _zz_10463;
  wire       [15:0]   _zz_10464;
  wire       [15:0]   _zz_10465;
  wire       [15:0]   _zz_10466;
  wire       [15:0]   _zz_10467;
  wire       [15:0]   _zz_10468;
  wire       [15:0]   _zz_10469;
  wire       [15:0]   _zz_10470;
  wire       [15:0]   _zz_10471;
  wire       [15:0]   _zz_10472;
  wire       [15:0]   _zz_10473;
  wire       [15:0]   _zz_10474;
  wire       [15:0]   _zz_10475;
  wire       [15:0]   _zz_10476;
  wire       [15:0]   _zz_10477;
  wire       [15:0]   _zz_10478;
  wire       [31:0]   _zz_10479;
  wire       [31:0]   _zz_10480;
  wire       [15:0]   _zz_10481;
  wire       [31:0]   _zz_10482;
  wire       [31:0]   _zz_10483;
  wire       [15:0]   _zz_10484;
  wire       [15:0]   _zz_10485;
  wire       [15:0]   _zz_10486;
  wire       [15:0]   _zz_10487;
  wire       [15:0]   _zz_10488;
  wire       [15:0]   _zz_10489;
  wire       [15:0]   _zz_10490;
  wire       [15:0]   _zz_10491;
  wire       [15:0]   _zz_10492;
  wire       [15:0]   _zz_10493;
  wire       [15:0]   _zz_10494;
  wire       [15:0]   _zz_10495;
  wire       [15:0]   _zz_10496;
  wire       [15:0]   _zz_10497;
  wire       [15:0]   _zz_10498;
  wire       [15:0]   _zz_10499;
  wire       [15:0]   _zz_10500;
  wire       [31:0]   _zz_10501;
  wire       [31:0]   _zz_10502;
  wire       [15:0]   _zz_10503;
  wire       [31:0]   _zz_10504;
  wire       [31:0]   _zz_10505;
  wire       [15:0]   _zz_10506;
  wire       [15:0]   _zz_10507;
  wire       [15:0]   _zz_10508;
  wire       [15:0]   _zz_10509;
  wire       [15:0]   _zz_10510;
  wire       [15:0]   _zz_10511;
  wire       [15:0]   _zz_10512;
  wire       [15:0]   _zz_10513;
  wire       [15:0]   _zz_10514;
  wire       [15:0]   _zz_10515;
  wire       [15:0]   _zz_10516;
  wire       [15:0]   _zz_10517;
  wire       [15:0]   _zz_10518;
  wire       [15:0]   _zz_10519;
  wire       [15:0]   _zz_10520;
  wire       [15:0]   _zz_10521;
  wire       [15:0]   _zz_10522;
  wire       [31:0]   _zz_10523;
  wire       [31:0]   _zz_10524;
  wire       [15:0]   _zz_10525;
  wire       [31:0]   _zz_10526;
  wire       [31:0]   _zz_10527;
  wire       [15:0]   _zz_10528;
  wire       [15:0]   _zz_10529;
  wire       [15:0]   _zz_10530;
  wire       [15:0]   _zz_10531;
  wire       [15:0]   _zz_10532;
  wire       [15:0]   _zz_10533;
  wire       [15:0]   _zz_10534;
  wire       [15:0]   _zz_10535;
  wire       [15:0]   _zz_10536;
  wire       [15:0]   _zz_10537;
  wire       [15:0]   _zz_10538;
  wire       [15:0]   _zz_10539;
  wire       [15:0]   _zz_10540;
  wire       [15:0]   _zz_10541;
  wire       [15:0]   _zz_10542;
  wire       [15:0]   _zz_10543;
  wire       [15:0]   _zz_10544;
  wire       [31:0]   _zz_10545;
  wire       [31:0]   _zz_10546;
  wire       [15:0]   _zz_10547;
  wire       [31:0]   _zz_10548;
  wire       [31:0]   _zz_10549;
  wire       [15:0]   _zz_10550;
  wire       [15:0]   _zz_10551;
  wire       [15:0]   _zz_10552;
  wire       [15:0]   _zz_10553;
  wire       [15:0]   _zz_10554;
  wire       [15:0]   _zz_10555;
  wire       [15:0]   _zz_10556;
  wire       [15:0]   _zz_10557;
  wire       [15:0]   _zz_10558;
  wire       [15:0]   _zz_10559;
  wire       [15:0]   _zz_10560;
  wire       [15:0]   _zz_10561;
  wire       [15:0]   _zz_10562;
  wire       [15:0]   _zz_10563;
  wire       [15:0]   _zz_10564;
  wire       [15:0]   _zz_10565;
  wire       [15:0]   _zz_10566;
  wire       [31:0]   _zz_10567;
  wire       [31:0]   _zz_10568;
  wire       [15:0]   _zz_10569;
  wire       [31:0]   _zz_10570;
  wire       [31:0]   _zz_10571;
  wire       [15:0]   _zz_10572;
  wire       [15:0]   _zz_10573;
  wire       [15:0]   _zz_10574;
  wire       [15:0]   _zz_10575;
  wire       [15:0]   _zz_10576;
  wire       [15:0]   _zz_10577;
  wire       [15:0]   _zz_10578;
  wire       [15:0]   _zz_10579;
  wire       [15:0]   _zz_10580;
  wire       [15:0]   _zz_10581;
  wire       [15:0]   _zz_10582;
  wire       [15:0]   _zz_10583;
  wire       [15:0]   _zz_10584;
  wire       [15:0]   _zz_10585;
  wire       [15:0]   _zz_10586;
  wire       [15:0]   _zz_10587;
  wire       [15:0]   _zz_10588;
  wire       [31:0]   _zz_10589;
  wire       [31:0]   _zz_10590;
  wire       [15:0]   _zz_10591;
  wire       [31:0]   _zz_10592;
  wire       [31:0]   _zz_10593;
  wire       [15:0]   _zz_10594;
  wire       [15:0]   _zz_10595;
  wire       [15:0]   _zz_10596;
  wire       [15:0]   _zz_10597;
  wire       [15:0]   _zz_10598;
  wire       [15:0]   _zz_10599;
  wire       [15:0]   _zz_10600;
  wire       [15:0]   _zz_10601;
  wire       [15:0]   _zz_10602;
  wire       [15:0]   _zz_10603;
  wire       [15:0]   _zz_10604;
  wire       [15:0]   _zz_10605;
  wire       [15:0]   _zz_10606;
  wire       [15:0]   _zz_10607;
  wire       [15:0]   _zz_10608;
  wire       [15:0]   _zz_10609;
  wire       [15:0]   _zz_10610;
  wire       [31:0]   _zz_10611;
  wire       [31:0]   _zz_10612;
  wire       [15:0]   _zz_10613;
  wire       [31:0]   _zz_10614;
  wire       [31:0]   _zz_10615;
  wire       [15:0]   _zz_10616;
  wire       [15:0]   _zz_10617;
  wire       [15:0]   _zz_10618;
  wire       [15:0]   _zz_10619;
  wire       [15:0]   _zz_10620;
  wire       [15:0]   _zz_10621;
  wire       [15:0]   _zz_10622;
  wire       [15:0]   _zz_10623;
  wire       [15:0]   _zz_10624;
  wire       [15:0]   _zz_10625;
  wire       [15:0]   _zz_10626;
  wire       [15:0]   _zz_10627;
  wire       [15:0]   _zz_10628;
  wire       [15:0]   _zz_10629;
  wire       [15:0]   _zz_10630;
  wire       [15:0]   _zz_10631;
  wire       [15:0]   _zz_10632;
  wire       [31:0]   _zz_10633;
  wire       [31:0]   _zz_10634;
  wire       [15:0]   _zz_10635;
  wire       [31:0]   _zz_10636;
  wire       [31:0]   _zz_10637;
  wire       [15:0]   _zz_10638;
  wire       [15:0]   _zz_10639;
  wire       [15:0]   _zz_10640;
  wire       [15:0]   _zz_10641;
  wire       [15:0]   _zz_10642;
  wire       [15:0]   _zz_10643;
  wire       [15:0]   _zz_10644;
  wire       [15:0]   _zz_10645;
  wire       [15:0]   _zz_10646;
  wire       [15:0]   _zz_10647;
  wire       [15:0]   _zz_10648;
  wire       [15:0]   _zz_10649;
  wire       [15:0]   _zz_10650;
  wire       [15:0]   _zz_10651;
  wire       [15:0]   _zz_10652;
  wire       [15:0]   _zz_10653;
  wire       [15:0]   _zz_10654;
  wire       [31:0]   _zz_10655;
  wire       [31:0]   _zz_10656;
  wire       [15:0]   _zz_10657;
  wire       [31:0]   _zz_10658;
  wire       [31:0]   _zz_10659;
  wire       [15:0]   _zz_10660;
  wire       [15:0]   _zz_10661;
  wire       [15:0]   _zz_10662;
  wire       [15:0]   _zz_10663;
  wire       [15:0]   _zz_10664;
  wire       [15:0]   _zz_10665;
  wire       [15:0]   _zz_10666;
  wire       [15:0]   _zz_10667;
  wire       [15:0]   _zz_10668;
  wire       [15:0]   _zz_10669;
  wire       [15:0]   _zz_10670;
  wire       [15:0]   _zz_10671;
  wire       [15:0]   _zz_10672;
  wire       [15:0]   _zz_10673;
  wire       [15:0]   _zz_10674;
  wire       [15:0]   _zz_10675;
  wire       [15:0]   _zz_10676;
  wire       [31:0]   _zz_10677;
  wire       [31:0]   _zz_10678;
  wire       [15:0]   _zz_10679;
  wire       [31:0]   _zz_10680;
  wire       [31:0]   _zz_10681;
  wire       [15:0]   _zz_10682;
  wire       [15:0]   _zz_10683;
  wire       [15:0]   _zz_10684;
  wire       [15:0]   _zz_10685;
  wire       [15:0]   _zz_10686;
  wire       [15:0]   _zz_10687;
  wire       [15:0]   _zz_10688;
  wire       [15:0]   _zz_10689;
  wire       [15:0]   _zz_10690;
  wire       [15:0]   _zz_10691;
  wire       [15:0]   _zz_10692;
  wire       [15:0]   _zz_10693;
  wire       [15:0]   _zz_10694;
  wire       [15:0]   _zz_10695;
  wire       [15:0]   _zz_10696;
  wire       [15:0]   _zz_10697;
  wire       [15:0]   _zz_10698;
  wire       [31:0]   _zz_10699;
  wire       [31:0]   _zz_10700;
  wire       [15:0]   _zz_10701;
  wire       [31:0]   _zz_10702;
  wire       [31:0]   _zz_10703;
  wire       [15:0]   _zz_10704;
  wire       [15:0]   _zz_10705;
  wire       [15:0]   _zz_10706;
  wire       [15:0]   _zz_10707;
  wire       [15:0]   _zz_10708;
  wire       [15:0]   _zz_10709;
  wire       [15:0]   _zz_10710;
  wire       [15:0]   _zz_10711;
  wire       [15:0]   _zz_10712;
  wire       [15:0]   _zz_10713;
  wire       [15:0]   _zz_10714;
  wire       [15:0]   _zz_10715;
  wire       [15:0]   _zz_10716;
  wire       [15:0]   _zz_10717;
  wire       [15:0]   _zz_10718;
  wire       [15:0]   _zz_10719;
  wire       [15:0]   _zz_10720;
  wire       [31:0]   _zz_10721;
  wire       [31:0]   _zz_10722;
  wire       [15:0]   _zz_10723;
  wire       [31:0]   _zz_10724;
  wire       [31:0]   _zz_10725;
  wire       [15:0]   _zz_10726;
  wire       [15:0]   _zz_10727;
  wire       [15:0]   _zz_10728;
  wire       [15:0]   _zz_10729;
  wire       [15:0]   _zz_10730;
  wire       [15:0]   _zz_10731;
  wire       [15:0]   _zz_10732;
  wire       [15:0]   _zz_10733;
  wire       [15:0]   _zz_10734;
  wire       [15:0]   _zz_10735;
  wire       [15:0]   _zz_10736;
  wire       [15:0]   _zz_10737;
  wire       [15:0]   _zz_10738;
  wire       [15:0]   _zz_10739;
  wire       [15:0]   _zz_10740;
  wire       [15:0]   _zz_10741;
  wire       [15:0]   _zz_10742;
  wire       [31:0]   _zz_10743;
  wire       [31:0]   _zz_10744;
  wire       [15:0]   _zz_10745;
  wire       [31:0]   _zz_10746;
  wire       [31:0]   _zz_10747;
  wire       [15:0]   _zz_10748;
  wire       [15:0]   _zz_10749;
  wire       [15:0]   _zz_10750;
  wire       [15:0]   _zz_10751;
  wire       [15:0]   _zz_10752;
  wire       [15:0]   _zz_10753;
  wire       [15:0]   _zz_10754;
  wire       [15:0]   _zz_10755;
  wire       [15:0]   _zz_10756;
  wire       [15:0]   _zz_10757;
  wire       [15:0]   _zz_10758;
  wire       [15:0]   _zz_10759;
  wire       [15:0]   _zz_10760;
  wire       [15:0]   _zz_10761;
  wire       [15:0]   _zz_10762;
  wire       [15:0]   _zz_10763;
  wire       [15:0]   _zz_10764;
  wire       [31:0]   _zz_10765;
  wire       [31:0]   _zz_10766;
  wire       [15:0]   _zz_10767;
  wire       [31:0]   _zz_10768;
  wire       [31:0]   _zz_10769;
  wire       [15:0]   _zz_10770;
  wire       [15:0]   _zz_10771;
  wire       [15:0]   _zz_10772;
  wire       [15:0]   _zz_10773;
  wire       [15:0]   _zz_10774;
  wire       [15:0]   _zz_10775;
  wire       [15:0]   _zz_10776;
  wire       [15:0]   _zz_10777;
  wire       [15:0]   _zz_10778;
  wire       [15:0]   _zz_10779;
  wire       [15:0]   _zz_10780;
  wire       [15:0]   _zz_10781;
  wire       [15:0]   _zz_10782;
  wire       [15:0]   _zz_10783;
  wire       [15:0]   _zz_10784;
  wire       [15:0]   _zz_10785;
  wire       [15:0]   _zz_10786;
  wire       [31:0]   _zz_10787;
  wire       [31:0]   _zz_10788;
  wire       [15:0]   _zz_10789;
  wire       [31:0]   _zz_10790;
  wire       [31:0]   _zz_10791;
  wire       [15:0]   _zz_10792;
  wire       [15:0]   _zz_10793;
  wire       [15:0]   _zz_10794;
  wire       [15:0]   _zz_10795;
  wire       [15:0]   _zz_10796;
  wire       [15:0]   _zz_10797;
  wire       [15:0]   _zz_10798;
  wire       [15:0]   _zz_10799;
  wire       [15:0]   _zz_10800;
  wire       [15:0]   _zz_10801;
  wire       [15:0]   _zz_10802;
  wire       [15:0]   _zz_10803;
  wire       [15:0]   _zz_10804;
  wire       [15:0]   _zz_10805;
  wire       [15:0]   _zz_10806;
  wire       [15:0]   _zz_10807;
  wire       [15:0]   _zz_10808;
  wire       [31:0]   _zz_10809;
  wire       [31:0]   _zz_10810;
  wire       [15:0]   _zz_10811;
  wire       [31:0]   _zz_10812;
  wire       [31:0]   _zz_10813;
  wire       [15:0]   _zz_10814;
  wire       [15:0]   _zz_10815;
  wire       [15:0]   _zz_10816;
  wire       [15:0]   _zz_10817;
  wire       [15:0]   _zz_10818;
  wire       [15:0]   _zz_10819;
  wire       [15:0]   _zz_10820;
  wire       [15:0]   _zz_10821;
  wire       [15:0]   _zz_10822;
  wire       [15:0]   _zz_10823;
  wire       [15:0]   _zz_10824;
  wire       [15:0]   _zz_10825;
  wire       [15:0]   _zz_10826;
  wire       [15:0]   _zz_10827;
  wire       [15:0]   _zz_10828;
  wire       [15:0]   _zz_10829;
  wire       [15:0]   _zz_10830;
  wire       [31:0]   _zz_10831;
  wire       [31:0]   _zz_10832;
  wire       [15:0]   _zz_10833;
  wire       [31:0]   _zz_10834;
  wire       [31:0]   _zz_10835;
  wire       [15:0]   _zz_10836;
  wire       [15:0]   _zz_10837;
  wire       [15:0]   _zz_10838;
  wire       [15:0]   _zz_10839;
  wire       [15:0]   _zz_10840;
  wire       [15:0]   _zz_10841;
  wire       [15:0]   _zz_10842;
  wire       [15:0]   _zz_10843;
  wire       [15:0]   _zz_10844;
  wire       [15:0]   _zz_10845;
  wire       [15:0]   _zz_10846;
  wire       [15:0]   _zz_10847;
  wire       [15:0]   _zz_10848;
  wire       [15:0]   _zz_10849;
  wire       [15:0]   _zz_10850;
  wire       [15:0]   _zz_10851;
  wire       [15:0]   _zz_10852;
  wire       [31:0]   _zz_10853;
  wire       [31:0]   _zz_10854;
  wire       [15:0]   _zz_10855;
  wire       [31:0]   _zz_10856;
  wire       [31:0]   _zz_10857;
  wire       [15:0]   _zz_10858;
  wire       [15:0]   _zz_10859;
  wire       [15:0]   _zz_10860;
  wire       [15:0]   _zz_10861;
  wire       [15:0]   _zz_10862;
  wire       [15:0]   _zz_10863;
  wire       [15:0]   _zz_10864;
  wire       [15:0]   _zz_10865;
  wire       [15:0]   _zz_10866;
  wire       [15:0]   _zz_10867;
  wire       [15:0]   _zz_10868;
  wire       [15:0]   _zz_10869;
  wire       [15:0]   _zz_10870;
  wire       [15:0]   _zz_10871;
  wire       [15:0]   _zz_10872;
  wire       [15:0]   _zz_10873;
  wire       [15:0]   _zz_10874;
  wire       [31:0]   _zz_10875;
  wire       [31:0]   _zz_10876;
  wire       [15:0]   _zz_10877;
  wire       [31:0]   _zz_10878;
  wire       [31:0]   _zz_10879;
  wire       [15:0]   _zz_10880;
  wire       [15:0]   _zz_10881;
  wire       [15:0]   _zz_10882;
  wire       [15:0]   _zz_10883;
  wire       [15:0]   _zz_10884;
  wire       [15:0]   _zz_10885;
  wire       [15:0]   _zz_10886;
  wire       [15:0]   _zz_10887;
  wire       [15:0]   _zz_10888;
  wire       [15:0]   _zz_10889;
  wire       [15:0]   _zz_10890;
  wire       [15:0]   _zz_10891;
  wire       [15:0]   _zz_10892;
  wire       [15:0]   _zz_10893;
  wire       [15:0]   _zz_10894;
  wire       [15:0]   _zz_10895;
  wire       [15:0]   _zz_10896;
  wire       [31:0]   _zz_10897;
  wire       [31:0]   _zz_10898;
  wire       [15:0]   _zz_10899;
  wire       [31:0]   _zz_10900;
  wire       [31:0]   _zz_10901;
  wire       [15:0]   _zz_10902;
  wire       [15:0]   _zz_10903;
  wire       [15:0]   _zz_10904;
  wire       [15:0]   _zz_10905;
  wire       [15:0]   _zz_10906;
  wire       [15:0]   _zz_10907;
  wire       [15:0]   _zz_10908;
  wire       [15:0]   _zz_10909;
  wire       [15:0]   _zz_10910;
  wire       [15:0]   _zz_10911;
  wire       [15:0]   _zz_10912;
  wire       [15:0]   _zz_10913;
  wire       [15:0]   _zz_10914;
  wire       [15:0]   _zz_10915;
  wire       [15:0]   _zz_10916;
  wire       [15:0]   _zz_10917;
  wire       [15:0]   _zz_10918;
  wire       [31:0]   _zz_10919;
  wire       [31:0]   _zz_10920;
  wire       [15:0]   _zz_10921;
  wire       [31:0]   _zz_10922;
  wire       [31:0]   _zz_10923;
  wire       [15:0]   _zz_10924;
  wire       [15:0]   _zz_10925;
  wire       [15:0]   _zz_10926;
  wire       [15:0]   _zz_10927;
  wire       [15:0]   _zz_10928;
  wire       [15:0]   _zz_10929;
  wire       [15:0]   _zz_10930;
  wire       [15:0]   _zz_10931;
  wire       [15:0]   _zz_10932;
  wire       [15:0]   _zz_10933;
  wire       [15:0]   _zz_10934;
  wire       [15:0]   _zz_10935;
  wire       [15:0]   _zz_10936;
  wire       [15:0]   _zz_10937;
  wire       [15:0]   _zz_10938;
  wire       [15:0]   _zz_10939;
  wire       [15:0]   _zz_10940;
  wire       [31:0]   _zz_10941;
  wire       [31:0]   _zz_10942;
  wire       [15:0]   _zz_10943;
  wire       [31:0]   _zz_10944;
  wire       [31:0]   _zz_10945;
  wire       [15:0]   _zz_10946;
  wire       [15:0]   _zz_10947;
  wire       [15:0]   _zz_10948;
  wire       [15:0]   _zz_10949;
  wire       [15:0]   _zz_10950;
  wire       [15:0]   _zz_10951;
  wire       [15:0]   _zz_10952;
  wire       [15:0]   _zz_10953;
  wire       [15:0]   _zz_10954;
  wire       [15:0]   _zz_10955;
  wire       [15:0]   _zz_10956;
  wire       [15:0]   _zz_10957;
  wire       [15:0]   _zz_10958;
  wire       [15:0]   _zz_10959;
  wire       [15:0]   _zz_10960;
  wire       [15:0]   _zz_10961;
  wire       [15:0]   _zz_10962;
  wire       [31:0]   _zz_10963;
  wire       [31:0]   _zz_10964;
  wire       [15:0]   _zz_10965;
  wire       [31:0]   _zz_10966;
  wire       [31:0]   _zz_10967;
  wire       [15:0]   _zz_10968;
  wire       [15:0]   _zz_10969;
  wire       [15:0]   _zz_10970;
  wire       [15:0]   _zz_10971;
  wire       [15:0]   _zz_10972;
  wire       [15:0]   _zz_10973;
  wire       [15:0]   _zz_10974;
  wire       [15:0]   _zz_10975;
  wire       [15:0]   _zz_10976;
  wire       [15:0]   _zz_10977;
  wire       [15:0]   _zz_10978;
  wire       [15:0]   _zz_10979;
  wire       [15:0]   _zz_10980;
  wire       [15:0]   _zz_10981;
  wire       [15:0]   _zz_10982;
  wire       [15:0]   _zz_10983;
  wire       [15:0]   _zz_10984;
  wire       [31:0]   _zz_10985;
  wire       [31:0]   _zz_10986;
  wire       [15:0]   _zz_10987;
  wire       [31:0]   _zz_10988;
  wire       [31:0]   _zz_10989;
  wire       [15:0]   _zz_10990;
  wire       [15:0]   _zz_10991;
  wire       [15:0]   _zz_10992;
  wire       [15:0]   _zz_10993;
  wire       [15:0]   _zz_10994;
  wire       [15:0]   _zz_10995;
  wire       [15:0]   _zz_10996;
  wire       [15:0]   _zz_10997;
  wire       [15:0]   _zz_10998;
  wire       [15:0]   _zz_10999;
  wire       [15:0]   _zz_11000;
  wire       [15:0]   _zz_11001;
  wire       [15:0]   _zz_11002;
  wire       [15:0]   _zz_11003;
  wire       [15:0]   _zz_11004;
  wire       [15:0]   _zz_11005;
  wire       [15:0]   _zz_11006;
  wire       [31:0]   _zz_11007;
  wire       [31:0]   _zz_11008;
  wire       [15:0]   _zz_11009;
  wire       [31:0]   _zz_11010;
  wire       [31:0]   _zz_11011;
  wire       [15:0]   _zz_11012;
  wire       [15:0]   _zz_11013;
  wire       [15:0]   _zz_11014;
  wire       [15:0]   _zz_11015;
  wire       [15:0]   _zz_11016;
  wire       [15:0]   _zz_11017;
  wire       [15:0]   _zz_11018;
  wire       [15:0]   _zz_11019;
  wire       [15:0]   _zz_11020;
  wire       [15:0]   _zz_11021;
  wire       [15:0]   _zz_11022;
  wire       [15:0]   _zz_11023;
  wire       [15:0]   _zz_11024;
  wire       [15:0]   _zz_11025;
  wire       [15:0]   _zz_11026;
  wire       [15:0]   _zz_11027;
  wire       [15:0]   _zz_11028;
  wire       [31:0]   _zz_11029;
  wire       [31:0]   _zz_11030;
  wire       [15:0]   _zz_11031;
  wire       [31:0]   _zz_11032;
  wire       [31:0]   _zz_11033;
  wire       [15:0]   _zz_11034;
  wire       [15:0]   _zz_11035;
  wire       [15:0]   _zz_11036;
  wire       [15:0]   _zz_11037;
  wire       [15:0]   _zz_11038;
  wire       [15:0]   _zz_11039;
  wire       [15:0]   _zz_11040;
  wire       [15:0]   _zz_11041;
  wire       [15:0]   _zz_11042;
  wire       [15:0]   _zz_11043;
  wire       [15:0]   _zz_11044;
  wire       [15:0]   _zz_11045;
  wire       [15:0]   _zz_11046;
  wire       [15:0]   _zz_11047;
  wire       [15:0]   _zz_11048;
  wire       [15:0]   _zz_11049;
  wire       [15:0]   _zz_11050;
  wire       [31:0]   _zz_11051;
  wire       [31:0]   _zz_11052;
  wire       [15:0]   _zz_11053;
  wire       [31:0]   _zz_11054;
  wire       [31:0]   _zz_11055;
  wire       [15:0]   _zz_11056;
  wire       [15:0]   _zz_11057;
  wire       [15:0]   _zz_11058;
  wire       [15:0]   _zz_11059;
  wire       [15:0]   _zz_11060;
  wire       [15:0]   _zz_11061;
  wire       [15:0]   _zz_11062;
  wire       [15:0]   _zz_11063;
  wire       [15:0]   _zz_11064;
  wire       [15:0]   _zz_11065;
  wire       [15:0]   _zz_11066;
  wire       [15:0]   _zz_11067;
  wire       [15:0]   _zz_11068;
  wire       [15:0]   _zz_11069;
  wire       [15:0]   _zz_11070;
  wire       [15:0]   _zz_11071;
  wire       [15:0]   _zz_11072;
  wire       [31:0]   _zz_11073;
  wire       [31:0]   _zz_11074;
  wire       [15:0]   _zz_11075;
  wire       [31:0]   _zz_11076;
  wire       [31:0]   _zz_11077;
  wire       [15:0]   _zz_11078;
  wire       [15:0]   _zz_11079;
  wire       [15:0]   _zz_11080;
  wire       [15:0]   _zz_11081;
  wire       [15:0]   _zz_11082;
  wire       [15:0]   _zz_11083;
  wire       [15:0]   _zz_11084;
  wire       [15:0]   _zz_11085;
  wire       [15:0]   _zz_11086;
  wire       [15:0]   _zz_11087;
  wire       [15:0]   _zz_11088;
  wire       [15:0]   _zz_11089;
  wire       [15:0]   _zz_11090;
  wire       [15:0]   _zz_11091;
  wire       [15:0]   _zz_11092;
  wire       [15:0]   _zz_11093;
  wire       [15:0]   _zz_11094;
  wire       [31:0]   _zz_11095;
  wire       [31:0]   _zz_11096;
  wire       [15:0]   _zz_11097;
  wire       [31:0]   _zz_11098;
  wire       [31:0]   _zz_11099;
  wire       [15:0]   _zz_11100;
  wire       [15:0]   _zz_11101;
  wire       [15:0]   _zz_11102;
  wire       [15:0]   _zz_11103;
  wire       [15:0]   _zz_11104;
  wire       [15:0]   _zz_11105;
  wire       [15:0]   _zz_11106;
  wire       [15:0]   _zz_11107;
  wire       [15:0]   _zz_11108;
  wire       [15:0]   _zz_11109;
  wire       [15:0]   _zz_11110;
  wire       [15:0]   _zz_11111;
  wire       [15:0]   _zz_11112;
  wire       [15:0]   _zz_11113;
  wire       [15:0]   _zz_11114;
  wire       [15:0]   _zz_11115;
  wire       [15:0]   _zz_11116;
  wire       [31:0]   _zz_11117;
  wire       [31:0]   _zz_11118;
  wire       [15:0]   _zz_11119;
  wire       [31:0]   _zz_11120;
  wire       [31:0]   _zz_11121;
  wire       [15:0]   _zz_11122;
  wire       [15:0]   _zz_11123;
  wire       [15:0]   _zz_11124;
  wire       [15:0]   _zz_11125;
  wire       [15:0]   _zz_11126;
  wire       [15:0]   _zz_11127;
  wire       [15:0]   _zz_11128;
  wire       [15:0]   _zz_11129;
  wire       [15:0]   _zz_11130;
  wire       [15:0]   _zz_11131;
  wire       [15:0]   _zz_11132;
  wire       [15:0]   _zz_11133;
  wire       [15:0]   _zz_11134;
  wire       [15:0]   _zz_11135;
  wire       [15:0]   _zz_11136;
  wire       [15:0]   _zz_11137;
  wire       [15:0]   _zz_11138;
  wire       [31:0]   _zz_11139;
  wire       [31:0]   _zz_11140;
  wire       [15:0]   _zz_11141;
  wire       [31:0]   _zz_11142;
  wire       [31:0]   _zz_11143;
  wire       [15:0]   _zz_11144;
  wire       [15:0]   _zz_11145;
  wire       [15:0]   _zz_11146;
  wire       [15:0]   _zz_11147;
  wire       [15:0]   _zz_11148;
  wire       [15:0]   _zz_11149;
  wire       [15:0]   _zz_11150;
  wire       [15:0]   _zz_11151;
  wire       [15:0]   _zz_11152;
  wire       [15:0]   _zz_11153;
  wire       [15:0]   _zz_11154;
  wire       [15:0]   _zz_11155;
  wire       [15:0]   _zz_11156;
  wire       [15:0]   _zz_11157;
  wire       [15:0]   _zz_11158;
  wire       [15:0]   _zz_11159;
  wire       [15:0]   _zz_11160;
  wire       [31:0]   _zz_11161;
  wire       [31:0]   _zz_11162;
  wire       [15:0]   _zz_11163;
  wire       [31:0]   _zz_11164;
  wire       [31:0]   _zz_11165;
  wire       [15:0]   _zz_11166;
  wire       [15:0]   _zz_11167;
  wire       [15:0]   _zz_11168;
  wire       [15:0]   _zz_11169;
  wire       [15:0]   _zz_11170;
  wire       [15:0]   _zz_11171;
  wire       [15:0]   _zz_11172;
  wire       [15:0]   _zz_11173;
  wire       [15:0]   _zz_11174;
  wire       [15:0]   _zz_11175;
  wire       [15:0]   _zz_11176;
  wire       [15:0]   _zz_11177;
  wire       [15:0]   _zz_11178;
  wire       [15:0]   _zz_11179;
  wire       [15:0]   _zz_11180;
  wire       [15:0]   _zz_11181;
  wire       [15:0]   _zz_11182;
  wire       [31:0]   _zz_11183;
  wire       [31:0]   _zz_11184;
  wire       [15:0]   _zz_11185;
  wire       [31:0]   _zz_11186;
  wire       [31:0]   _zz_11187;
  wire       [15:0]   _zz_11188;
  wire       [15:0]   _zz_11189;
  wire       [15:0]   _zz_11190;
  wire       [15:0]   _zz_11191;
  wire       [15:0]   _zz_11192;
  wire       [15:0]   _zz_11193;
  wire       [15:0]   _zz_11194;
  wire       [15:0]   _zz_11195;
  wire       [15:0]   _zz_11196;
  wire       [15:0]   _zz_11197;
  wire       [15:0]   _zz_11198;
  wire       [15:0]   _zz_11199;
  wire       [15:0]   _zz_11200;
  wire       [15:0]   _zz_11201;
  wire       [15:0]   _zz_11202;
  wire       [15:0]   _zz_11203;
  wire       [15:0]   _zz_11204;
  wire       [31:0]   _zz_11205;
  wire       [31:0]   _zz_11206;
  wire       [15:0]   _zz_11207;
  wire       [31:0]   _zz_11208;
  wire       [31:0]   _zz_11209;
  wire       [15:0]   _zz_11210;
  wire       [15:0]   _zz_11211;
  wire       [15:0]   _zz_11212;
  wire       [15:0]   _zz_11213;
  wire       [15:0]   _zz_11214;
  wire       [15:0]   _zz_11215;
  wire       [15:0]   _zz_11216;
  wire       [15:0]   _zz_11217;
  wire       [15:0]   _zz_11218;
  wire       [15:0]   _zz_11219;
  wire       [15:0]   _zz_11220;
  wire       [15:0]   _zz_11221;
  wire       [15:0]   _zz_11222;
  wire       [15:0]   _zz_11223;
  wire       [15:0]   _zz_11224;
  wire       [15:0]   _zz_11225;
  wire       [15:0]   _zz_11226;
  wire       [31:0]   _zz_11227;
  wire       [31:0]   _zz_11228;
  wire       [15:0]   _zz_11229;
  wire       [31:0]   _zz_11230;
  wire       [31:0]   _zz_11231;
  wire       [15:0]   _zz_11232;
  wire       [15:0]   _zz_11233;
  wire       [15:0]   _zz_11234;
  wire       [15:0]   _zz_11235;
  wire       [15:0]   _zz_11236;
  wire       [15:0]   _zz_11237;
  wire       [15:0]   _zz_11238;
  wire       [15:0]   _zz_11239;
  wire       [15:0]   _zz_11240;
  wire       [15:0]   _zz_11241;
  wire       [15:0]   _zz_11242;
  wire       [15:0]   _zz_11243;
  wire       [15:0]   _zz_11244;
  wire       [15:0]   _zz_11245;
  wire       [15:0]   _zz_11246;
  wire       [15:0]   _zz_11247;
  wire       [15:0]   _zz_11248;
  wire       [31:0]   _zz_11249;
  wire       [31:0]   _zz_11250;
  wire       [15:0]   _zz_11251;
  wire       [31:0]   _zz_11252;
  wire       [31:0]   _zz_11253;
  wire       [15:0]   _zz_11254;
  wire       [15:0]   _zz_11255;
  wire       [15:0]   _zz_11256;
  wire       [15:0]   _zz_11257;
  wire       [15:0]   _zz_11258;
  wire       [15:0]   _zz_11259;
  wire       [15:0]   _zz_11260;
  wire       [15:0]   _zz_11261;
  wire       [15:0]   _zz_11262;
  wire       [15:0]   _zz_11263;
  wire       [15:0]   _zz_11264;
  wire       [15:0]   _zz_11265;
  wire       [15:0]   _zz_11266;
  wire       [15:0]   _zz_11267;
  wire       [15:0]   _zz_11268;
  wire       [15:0]   _zz_11269;
  wire       [15:0]   _zz_11270;
  wire       [31:0]   _zz_11271;
  wire       [31:0]   _zz_11272;
  wire       [15:0]   _zz_11273;
  wire       [31:0]   _zz_11274;
  wire       [31:0]   _zz_11275;
  wire       [15:0]   _zz_11276;
  wire       [15:0]   _zz_11277;
  wire       [15:0]   _zz_11278;
  wire       [15:0]   _zz_11279;
  wire       [15:0]   _zz_11280;
  wire       [15:0]   _zz_11281;
  wire       [15:0]   _zz_11282;
  wire       [15:0]   _zz_11283;
  wire       [15:0]   _zz_11284;
  wire       [15:0]   _zz_11285;
  wire       [15:0]   _zz_11286;
  wire       [15:0]   _zz_11287;
  wire       [15:0]   _zz_11288;
  wire       [15:0]   _zz_11289;
  wire       [15:0]   _zz_11290;
  wire       [15:0]   _zz_11291;
  wire       [15:0]   _zz_11292;
  wire       [31:0]   _zz_11293;
  wire       [31:0]   _zz_11294;
  wire       [15:0]   _zz_11295;
  wire       [31:0]   _zz_11296;
  wire       [31:0]   _zz_11297;
  wire       [15:0]   _zz_11298;
  wire       [15:0]   _zz_11299;
  wire       [15:0]   _zz_11300;
  wire       [15:0]   _zz_11301;
  wire       [15:0]   _zz_11302;
  wire       [15:0]   _zz_11303;
  wire       [15:0]   _zz_11304;
  wire       [15:0]   _zz_11305;
  wire       [15:0]   _zz_11306;
  wire       [15:0]   _zz_11307;
  wire       [15:0]   _zz_11308;
  wire       [15:0]   _zz_11309;
  wire       [15:0]   _zz_11310;
  wire       [15:0]   _zz_11311;
  wire       [15:0]   _zz_11312;
  wire       [15:0]   _zz_11313;
  wire       [15:0]   _zz_11314;
  wire       [31:0]   _zz_11315;
  wire       [31:0]   _zz_11316;
  wire       [15:0]   _zz_11317;
  wire       [31:0]   _zz_11318;
  wire       [31:0]   _zz_11319;
  wire       [15:0]   _zz_11320;
  wire       [15:0]   _zz_11321;
  wire       [15:0]   _zz_11322;
  wire       [15:0]   _zz_11323;
  wire       [15:0]   _zz_11324;
  wire       [15:0]   _zz_11325;
  wire       [15:0]   _zz_11326;
  wire       [15:0]   _zz_11327;
  wire       [15:0]   _zz_11328;
  wire       [15:0]   _zz_11329;
  wire       [15:0]   _zz_11330;
  wire       [15:0]   _zz_11331;
  wire       [15:0]   _zz_11332;
  wire       [15:0]   _zz_11333;
  wire       [15:0]   _zz_11334;
  wire       [15:0]   _zz_11335;
  wire       [15:0]   _zz_11336;
  wire       [31:0]   _zz_11337;
  wire       [31:0]   _zz_11338;
  wire       [15:0]   _zz_11339;
  wire       [31:0]   _zz_11340;
  wire       [31:0]   _zz_11341;
  wire       [15:0]   _zz_11342;
  wire       [15:0]   _zz_11343;
  wire       [15:0]   _zz_11344;
  wire       [15:0]   _zz_11345;
  wire       [15:0]   _zz_11346;
  wire       [15:0]   _zz_11347;
  wire       [15:0]   _zz_11348;
  wire       [15:0]   _zz_11349;
  wire       [15:0]   _zz_11350;
  wire       [15:0]   _zz_11351;
  wire       [15:0]   _zz_11352;
  wire       [15:0]   _zz_11353;
  wire       [15:0]   _zz_11354;
  wire       [15:0]   _zz_11355;
  wire       [15:0]   _zz_11356;
  wire       [15:0]   _zz_11357;
  wire       [15:0]   _zz_11358;
  wire       [31:0]   _zz_11359;
  wire       [31:0]   _zz_11360;
  wire       [15:0]   _zz_11361;
  wire       [31:0]   _zz_11362;
  wire       [31:0]   _zz_11363;
  wire       [15:0]   _zz_11364;
  wire       [15:0]   _zz_11365;
  wire       [15:0]   _zz_11366;
  wire       [15:0]   _zz_11367;
  wire       [15:0]   _zz_11368;
  wire       [15:0]   _zz_11369;
  wire       [15:0]   _zz_11370;
  wire       [15:0]   _zz_11371;
  wire       [15:0]   _zz_11372;
  wire       [15:0]   _zz_11373;
  wire       [15:0]   _zz_11374;
  wire       [15:0]   _zz_11375;
  wire       [15:0]   _zz_11376;
  wire       [15:0]   _zz_11377;
  wire       [15:0]   _zz_11378;
  wire       [15:0]   _zz_11379;
  wire       [15:0]   _zz_11380;
  wire       [31:0]   _zz_11381;
  wire       [31:0]   _zz_11382;
  wire       [15:0]   _zz_11383;
  wire       [31:0]   _zz_11384;
  wire       [31:0]   _zz_11385;
  wire       [15:0]   _zz_11386;
  wire       [15:0]   _zz_11387;
  wire       [15:0]   _zz_11388;
  wire       [15:0]   _zz_11389;
  wire       [15:0]   _zz_11390;
  wire       [15:0]   _zz_11391;
  wire       [15:0]   _zz_11392;
  wire       [15:0]   _zz_11393;
  wire       [15:0]   _zz_11394;
  wire       [15:0]   _zz_11395;
  wire       [15:0]   _zz_11396;
  wire       [15:0]   _zz_11397;
  wire       [15:0]   _zz_11398;
  wire       [15:0]   _zz_11399;
  wire       [15:0]   _zz_11400;
  wire       [15:0]   _zz_11401;
  wire       [15:0]   _zz_11402;
  wire       [31:0]   _zz_11403;
  wire       [31:0]   _zz_11404;
  wire       [15:0]   _zz_11405;
  wire       [31:0]   _zz_11406;
  wire       [31:0]   _zz_11407;
  wire       [15:0]   _zz_11408;
  wire       [15:0]   _zz_11409;
  wire       [15:0]   _zz_11410;
  wire       [15:0]   _zz_11411;
  wire       [15:0]   _zz_11412;
  wire       [15:0]   _zz_11413;
  wire       [15:0]   _zz_11414;
  wire       [15:0]   _zz_11415;
  wire       [15:0]   _zz_11416;
  wire       [15:0]   _zz_11417;
  wire       [15:0]   _zz_11418;
  wire       [15:0]   _zz_11419;
  wire       [15:0]   _zz_11420;
  wire       [15:0]   _zz_11421;
  wire       [15:0]   _zz_11422;
  wire       [15:0]   _zz_11423;
  wire       [15:0]   _zz_11424;
  wire       [31:0]   _zz_11425;
  wire       [31:0]   _zz_11426;
  wire       [15:0]   _zz_11427;
  wire       [31:0]   _zz_11428;
  wire       [31:0]   _zz_11429;
  wire       [15:0]   _zz_11430;
  wire       [15:0]   _zz_11431;
  wire       [15:0]   _zz_11432;
  wire       [15:0]   _zz_11433;
  wire       [15:0]   _zz_11434;
  wire       [15:0]   _zz_11435;
  wire       [15:0]   _zz_11436;
  wire       [15:0]   _zz_11437;
  wire       [15:0]   _zz_11438;
  wire       [15:0]   _zz_11439;
  wire       [15:0]   _zz_11440;
  wire       [15:0]   _zz_11441;
  wire       [15:0]   _zz_11442;
  wire       [15:0]   _zz_11443;
  wire       [15:0]   _zz_11444;
  wire       [15:0]   _zz_11445;
  wire       [15:0]   _zz_11446;
  wire       [31:0]   _zz_11447;
  wire       [31:0]   _zz_11448;
  wire       [15:0]   _zz_11449;
  wire       [31:0]   _zz_11450;
  wire       [31:0]   _zz_11451;
  wire       [15:0]   _zz_11452;
  wire       [15:0]   _zz_11453;
  wire       [15:0]   _zz_11454;
  wire       [15:0]   _zz_11455;
  wire       [15:0]   _zz_11456;
  wire       [15:0]   _zz_11457;
  wire       [15:0]   _zz_11458;
  wire       [15:0]   _zz_11459;
  wire       [15:0]   _zz_11460;
  wire       [15:0]   _zz_11461;
  wire       [15:0]   _zz_11462;
  wire       [15:0]   _zz_11463;
  wire       [15:0]   _zz_11464;
  wire       [15:0]   _zz_11465;
  wire       [15:0]   _zz_11466;
  wire       [15:0]   _zz_11467;
  wire       [15:0]   _zz_11468;
  wire       [31:0]   _zz_11469;
  wire       [31:0]   _zz_11470;
  wire       [15:0]   _zz_11471;
  wire       [31:0]   _zz_11472;
  wire       [31:0]   _zz_11473;
  wire       [15:0]   _zz_11474;
  wire       [15:0]   _zz_11475;
  wire       [15:0]   _zz_11476;
  wire       [15:0]   _zz_11477;
  wire       [15:0]   _zz_11478;
  wire       [15:0]   _zz_11479;
  wire       [15:0]   _zz_11480;
  wire       [15:0]   _zz_11481;
  wire       [15:0]   _zz_11482;
  wire       [15:0]   _zz_11483;
  wire       [15:0]   _zz_11484;
  wire       [15:0]   _zz_11485;
  wire       [15:0]   _zz_11486;
  wire       [15:0]   _zz_11487;
  wire       [15:0]   _zz_11488;
  wire       [15:0]   _zz_11489;
  wire       [15:0]   _zz_11490;
  wire       [31:0]   _zz_11491;
  wire       [31:0]   _zz_11492;
  wire       [15:0]   _zz_11493;
  wire       [31:0]   _zz_11494;
  wire       [31:0]   _zz_11495;
  wire       [15:0]   _zz_11496;
  wire       [15:0]   _zz_11497;
  wire       [15:0]   _zz_11498;
  wire       [15:0]   _zz_11499;
  wire       [15:0]   _zz_11500;
  wire       [15:0]   _zz_11501;
  wire       [15:0]   _zz_11502;
  wire       [15:0]   _zz_11503;
  wire       [15:0]   _zz_11504;
  wire       [15:0]   _zz_11505;
  wire       [15:0]   _zz_11506;
  wire       [15:0]   _zz_11507;
  wire       [15:0]   _zz_11508;
  wire       [15:0]   _zz_11509;
  wire       [15:0]   _zz_11510;
  wire       [15:0]   _zz_11511;
  wire       [15:0]   _zz_11512;
  wire       [31:0]   _zz_11513;
  wire       [31:0]   _zz_11514;
  wire       [15:0]   _zz_11515;
  wire       [31:0]   _zz_11516;
  wire       [31:0]   _zz_11517;
  wire       [15:0]   _zz_11518;
  wire       [15:0]   _zz_11519;
  wire       [15:0]   _zz_11520;
  wire       [15:0]   _zz_11521;
  wire       [15:0]   _zz_11522;
  wire       [15:0]   _zz_11523;
  wire       [15:0]   _zz_11524;
  wire       [15:0]   _zz_11525;
  wire       [15:0]   _zz_11526;
  wire       [15:0]   _zz_11527;
  wire       [15:0]   _zz_11528;
  wire       [15:0]   _zz_11529;
  wire       [15:0]   _zz_11530;
  wire       [15:0]   _zz_11531;
  wire       [15:0]   _zz_11532;
  wire       [15:0]   _zz_11533;
  wire       [15:0]   _zz_11534;
  wire       [31:0]   _zz_11535;
  wire       [31:0]   _zz_11536;
  wire       [15:0]   _zz_11537;
  wire       [31:0]   _zz_11538;
  wire       [31:0]   _zz_11539;
  wire       [15:0]   _zz_11540;
  wire       [15:0]   _zz_11541;
  wire       [15:0]   _zz_11542;
  wire       [15:0]   _zz_11543;
  wire       [15:0]   _zz_11544;
  wire       [15:0]   _zz_11545;
  wire       [15:0]   _zz_11546;
  wire       [15:0]   _zz_11547;
  wire       [15:0]   _zz_11548;
  wire       [15:0]   _zz_11549;
  wire       [15:0]   _zz_11550;
  wire       [15:0]   _zz_11551;
  wire       [15:0]   _zz_11552;
  wire       [15:0]   _zz_11553;
  wire       [15:0]   _zz_11554;
  wire       [15:0]   _zz_11555;
  wire       [15:0]   _zz_11556;
  wire       [31:0]   _zz_11557;
  wire       [31:0]   _zz_11558;
  wire       [15:0]   _zz_11559;
  wire       [31:0]   _zz_11560;
  wire       [31:0]   _zz_11561;
  wire       [15:0]   _zz_11562;
  wire       [15:0]   _zz_11563;
  wire       [15:0]   _zz_11564;
  wire       [15:0]   _zz_11565;
  wire       [15:0]   _zz_11566;
  wire       [15:0]   _zz_11567;
  wire       [15:0]   _zz_11568;
  wire       [15:0]   _zz_11569;
  wire       [15:0]   _zz_11570;
  wire       [15:0]   _zz_11571;
  wire       [15:0]   _zz_11572;
  wire       [15:0]   _zz_11573;
  wire       [15:0]   _zz_11574;
  wire       [15:0]   _zz_11575;
  wire       [15:0]   _zz_11576;
  wire       [15:0]   _zz_11577;
  wire       [15:0]   _zz_11578;
  wire       [31:0]   _zz_11579;
  wire       [31:0]   _zz_11580;
  wire       [15:0]   _zz_11581;
  wire       [31:0]   _zz_11582;
  wire       [31:0]   _zz_11583;
  wire       [15:0]   _zz_11584;
  wire       [15:0]   _zz_11585;
  wire       [15:0]   _zz_11586;
  wire       [15:0]   _zz_11587;
  wire       [15:0]   _zz_11588;
  wire       [15:0]   _zz_11589;
  wire       [15:0]   _zz_11590;
  wire       [15:0]   _zz_11591;
  wire       [15:0]   _zz_11592;
  wire       [15:0]   _zz_11593;
  wire       [15:0]   _zz_11594;
  wire       [15:0]   _zz_11595;
  wire       [15:0]   _zz_11596;
  wire       [15:0]   _zz_11597;
  wire       [15:0]   _zz_11598;
  wire       [15:0]   _zz_11599;
  wire       [15:0]   _zz_11600;
  wire       [31:0]   _zz_11601;
  wire       [31:0]   _zz_11602;
  wire       [15:0]   _zz_11603;
  wire       [31:0]   _zz_11604;
  wire       [31:0]   _zz_11605;
  wire       [15:0]   _zz_11606;
  wire       [15:0]   _zz_11607;
  wire       [15:0]   _zz_11608;
  wire       [15:0]   _zz_11609;
  wire       [15:0]   _zz_11610;
  wire       [15:0]   _zz_11611;
  wire       [15:0]   _zz_11612;
  wire       [15:0]   _zz_11613;
  wire       [15:0]   _zz_11614;
  wire       [15:0]   _zz_11615;
  wire       [15:0]   _zz_11616;
  wire       [15:0]   _zz_11617;
  wire       [15:0]   _zz_11618;
  wire       [15:0]   _zz_11619;
  wire       [15:0]   _zz_11620;
  wire       [15:0]   _zz_11621;
  wire       [15:0]   _zz_11622;
  wire       [31:0]   _zz_11623;
  wire       [31:0]   _zz_11624;
  wire       [15:0]   _zz_11625;
  wire       [31:0]   _zz_11626;
  wire       [31:0]   _zz_11627;
  wire       [15:0]   _zz_11628;
  wire       [15:0]   _zz_11629;
  wire       [15:0]   _zz_11630;
  wire       [15:0]   _zz_11631;
  wire       [15:0]   _zz_11632;
  wire       [15:0]   _zz_11633;
  wire       [15:0]   _zz_11634;
  wire       [15:0]   _zz_11635;
  wire       [15:0]   _zz_11636;
  wire       [15:0]   _zz_11637;
  wire       [15:0]   _zz_11638;
  wire       [15:0]   _zz_11639;
  wire       [15:0]   _zz_11640;
  wire       [15:0]   _zz_11641;
  wire       [15:0]   _zz_11642;
  wire       [15:0]   _zz_11643;
  wire       [15:0]   _zz_11644;
  wire       [31:0]   _zz_11645;
  wire       [31:0]   _zz_11646;
  wire       [15:0]   _zz_11647;
  wire       [31:0]   _zz_11648;
  wire       [31:0]   _zz_11649;
  wire       [15:0]   _zz_11650;
  wire       [15:0]   _zz_11651;
  wire       [15:0]   _zz_11652;
  wire       [15:0]   _zz_11653;
  wire       [15:0]   _zz_11654;
  wire       [15:0]   _zz_11655;
  wire       [15:0]   _zz_11656;
  wire       [15:0]   _zz_11657;
  wire       [15:0]   _zz_11658;
  wire       [15:0]   _zz_11659;
  wire       [15:0]   _zz_11660;
  wire       [15:0]   _zz_11661;
  wire       [15:0]   _zz_11662;
  wire       [15:0]   _zz_11663;
  wire       [15:0]   _zz_11664;
  wire       [15:0]   _zz_11665;
  wire       [15:0]   _zz_11666;
  wire       [31:0]   _zz_11667;
  wire       [31:0]   _zz_11668;
  wire       [15:0]   _zz_11669;
  wire       [31:0]   _zz_11670;
  wire       [31:0]   _zz_11671;
  wire       [15:0]   _zz_11672;
  wire       [15:0]   _zz_11673;
  wire       [15:0]   _zz_11674;
  wire       [15:0]   _zz_11675;
  wire       [15:0]   _zz_11676;
  wire       [15:0]   _zz_11677;
  wire       [15:0]   _zz_11678;
  wire       [15:0]   _zz_11679;
  wire       [15:0]   _zz_11680;
  wire       [15:0]   _zz_11681;
  wire       [15:0]   _zz_11682;
  wire       [15:0]   _zz_11683;
  wire       [15:0]   _zz_11684;
  wire       [15:0]   _zz_11685;
  wire       [15:0]   _zz_11686;
  wire       [15:0]   _zz_11687;
  wire       [15:0]   _zz_11688;
  wire       [31:0]   _zz_11689;
  wire       [31:0]   _zz_11690;
  wire       [15:0]   _zz_11691;
  wire       [31:0]   _zz_11692;
  wire       [31:0]   _zz_11693;
  wire       [15:0]   _zz_11694;
  wire       [15:0]   _zz_11695;
  wire       [15:0]   _zz_11696;
  wire       [15:0]   _zz_11697;
  wire       [15:0]   _zz_11698;
  wire       [15:0]   _zz_11699;
  wire       [15:0]   _zz_11700;
  wire       [15:0]   _zz_11701;
  wire       [15:0]   _zz_11702;
  wire       [15:0]   _zz_11703;
  wire       [15:0]   _zz_11704;
  wire       [15:0]   _zz_11705;
  wire       [15:0]   _zz_11706;
  wire       [15:0]   _zz_11707;
  wire       [15:0]   _zz_11708;
  wire       [15:0]   _zz_11709;
  wire       [15:0]   _zz_11710;
  wire       [31:0]   _zz_11711;
  wire       [31:0]   _zz_11712;
  wire       [15:0]   _zz_11713;
  wire       [31:0]   _zz_11714;
  wire       [31:0]   _zz_11715;
  wire       [15:0]   _zz_11716;
  wire       [15:0]   _zz_11717;
  wire       [15:0]   _zz_11718;
  wire       [15:0]   _zz_11719;
  wire       [15:0]   _zz_11720;
  wire       [15:0]   _zz_11721;
  wire       [15:0]   _zz_11722;
  wire       [15:0]   _zz_11723;
  wire       [15:0]   _zz_11724;
  wire       [15:0]   _zz_11725;
  wire       [15:0]   _zz_11726;
  wire       [15:0]   _zz_11727;
  wire       [15:0]   _zz_11728;
  wire       [15:0]   _zz_11729;
  wire       [15:0]   _zz_11730;
  wire       [15:0]   _zz_11731;
  wire       [15:0]   _zz_11732;
  wire       [31:0]   _zz_11733;
  wire       [31:0]   _zz_11734;
  wire       [15:0]   _zz_11735;
  wire       [31:0]   _zz_11736;
  wire       [31:0]   _zz_11737;
  wire       [15:0]   _zz_11738;
  wire       [15:0]   _zz_11739;
  wire       [15:0]   _zz_11740;
  wire       [15:0]   _zz_11741;
  wire       [15:0]   _zz_11742;
  wire       [15:0]   _zz_11743;
  wire       [15:0]   _zz_11744;
  wire       [15:0]   _zz_11745;
  wire       [15:0]   _zz_11746;
  wire       [15:0]   _zz_11747;
  wire       [15:0]   _zz_11748;
  wire       [15:0]   _zz_11749;
  wire       [15:0]   _zz_11750;
  wire       [15:0]   _zz_11751;
  wire       [15:0]   _zz_11752;
  wire       [15:0]   _zz_11753;
  wire       [15:0]   _zz_11754;
  wire       [31:0]   _zz_11755;
  wire       [31:0]   _zz_11756;
  wire       [15:0]   _zz_11757;
  wire       [31:0]   _zz_11758;
  wire       [31:0]   _zz_11759;
  wire       [15:0]   _zz_11760;
  wire       [15:0]   _zz_11761;
  wire       [15:0]   _zz_11762;
  wire       [15:0]   _zz_11763;
  wire       [15:0]   _zz_11764;
  wire       [15:0]   _zz_11765;
  wire       [15:0]   _zz_11766;
  wire       [15:0]   _zz_11767;
  wire       [15:0]   _zz_11768;
  wire       [15:0]   _zz_11769;
  wire       [15:0]   _zz_11770;
  wire       [15:0]   _zz_11771;
  wire       [15:0]   _zz_11772;
  wire       [15:0]   _zz_11773;
  wire       [15:0]   _zz_11774;
  wire       [15:0]   _zz_11775;
  wire       [15:0]   _zz_11776;
  wire       [31:0]   _zz_11777;
  wire       [31:0]   _zz_11778;
  wire       [15:0]   _zz_11779;
  wire       [31:0]   _zz_11780;
  wire       [31:0]   _zz_11781;
  wire       [15:0]   _zz_11782;
  wire       [15:0]   _zz_11783;
  wire       [15:0]   _zz_11784;
  wire       [15:0]   _zz_11785;
  wire       [15:0]   _zz_11786;
  wire       [15:0]   _zz_11787;
  wire       [15:0]   _zz_11788;
  wire       [15:0]   _zz_11789;
  wire       [15:0]   _zz_11790;
  wire       [15:0]   _zz_11791;
  wire       [15:0]   _zz_11792;
  wire       [15:0]   _zz_11793;
  wire       [15:0]   _zz_11794;
  wire       [15:0]   _zz_11795;
  wire       [15:0]   _zz_11796;
  wire       [15:0]   _zz_11797;
  wire       [15:0]   _zz_11798;
  wire       [31:0]   _zz_11799;
  wire       [31:0]   _zz_11800;
  wire       [15:0]   _zz_11801;
  wire       [31:0]   _zz_11802;
  wire       [31:0]   _zz_11803;
  wire       [15:0]   _zz_11804;
  wire       [15:0]   _zz_11805;
  wire       [15:0]   _zz_11806;
  wire       [15:0]   _zz_11807;
  wire       [15:0]   _zz_11808;
  wire       [15:0]   _zz_11809;
  wire       [15:0]   _zz_11810;
  wire       [15:0]   _zz_11811;
  wire       [15:0]   _zz_11812;
  wire       [15:0]   _zz_11813;
  wire       [15:0]   _zz_11814;
  wire       [15:0]   _zz_11815;
  wire       [15:0]   _zz_11816;
  wire       [15:0]   _zz_11817;
  wire       [15:0]   _zz_11818;
  wire       [15:0]   _zz_11819;
  wire       [15:0]   _zz_11820;
  wire       [31:0]   _zz_11821;
  wire       [31:0]   _zz_11822;
  wire       [15:0]   _zz_11823;
  wire       [31:0]   _zz_11824;
  wire       [31:0]   _zz_11825;
  wire       [15:0]   _zz_11826;
  wire       [15:0]   _zz_11827;
  wire       [15:0]   _zz_11828;
  wire       [15:0]   _zz_11829;
  wire       [15:0]   _zz_11830;
  wire       [15:0]   _zz_11831;
  wire       [15:0]   _zz_11832;
  wire       [15:0]   _zz_11833;
  wire       [15:0]   _zz_11834;
  wire       [15:0]   _zz_11835;
  wire       [15:0]   _zz_11836;
  wire       [15:0]   _zz_11837;
  wire       [15:0]   _zz_11838;
  wire       [15:0]   _zz_11839;
  wire       [15:0]   _zz_11840;
  wire       [15:0]   _zz_11841;
  wire       [15:0]   _zz_11842;
  wire       [31:0]   _zz_11843;
  wire       [31:0]   _zz_11844;
  wire       [15:0]   _zz_11845;
  wire       [31:0]   _zz_11846;
  wire       [31:0]   _zz_11847;
  wire       [15:0]   _zz_11848;
  wire       [15:0]   _zz_11849;
  wire       [15:0]   _zz_11850;
  wire       [15:0]   _zz_11851;
  wire       [15:0]   _zz_11852;
  wire       [15:0]   _zz_11853;
  wire       [15:0]   _zz_11854;
  wire       [15:0]   _zz_11855;
  wire       [15:0]   _zz_11856;
  wire       [15:0]   _zz_11857;
  wire       [15:0]   _zz_11858;
  wire       [15:0]   _zz_11859;
  wire       [15:0]   _zz_11860;
  wire       [15:0]   _zz_11861;
  wire       [15:0]   _zz_11862;
  wire       [15:0]   _zz_11863;
  wire       [15:0]   _zz_11864;
  wire       [31:0]   _zz_11865;
  wire       [31:0]   _zz_11866;
  wire       [15:0]   _zz_11867;
  wire       [31:0]   _zz_11868;
  wire       [31:0]   _zz_11869;
  wire       [15:0]   _zz_11870;
  wire       [15:0]   _zz_11871;
  wire       [15:0]   _zz_11872;
  wire       [15:0]   _zz_11873;
  wire       [15:0]   _zz_11874;
  wire       [15:0]   _zz_11875;
  wire       [15:0]   _zz_11876;
  wire       [15:0]   _zz_11877;
  wire       [15:0]   _zz_11878;
  wire       [15:0]   _zz_11879;
  wire       [15:0]   _zz_11880;
  wire       [15:0]   _zz_11881;
  wire       [15:0]   _zz_11882;
  wire       [15:0]   _zz_11883;
  wire       [15:0]   _zz_11884;
  wire       [15:0]   _zz_11885;
  wire       [15:0]   _zz_11886;
  wire       [31:0]   _zz_11887;
  wire       [31:0]   _zz_11888;
  wire       [15:0]   _zz_11889;
  wire       [31:0]   _zz_11890;
  wire       [31:0]   _zz_11891;
  wire       [15:0]   _zz_11892;
  wire       [15:0]   _zz_11893;
  wire       [15:0]   _zz_11894;
  wire       [15:0]   _zz_11895;
  wire       [15:0]   _zz_11896;
  wire       [15:0]   _zz_11897;
  wire       [15:0]   _zz_11898;
  wire       [15:0]   _zz_11899;
  wire       [15:0]   _zz_11900;
  wire       [15:0]   _zz_11901;
  wire       [15:0]   _zz_11902;
  wire       [15:0]   _zz_11903;
  wire       [15:0]   _zz_11904;
  wire       [15:0]   _zz_11905;
  wire       [15:0]   _zz_11906;
  wire       [15:0]   _zz_11907;
  wire       [15:0]   _zz_11908;
  wire       [31:0]   _zz_11909;
  wire       [31:0]   _zz_11910;
  wire       [15:0]   _zz_11911;
  wire       [31:0]   _zz_11912;
  wire       [31:0]   _zz_11913;
  wire       [15:0]   _zz_11914;
  wire       [15:0]   _zz_11915;
  wire       [15:0]   _zz_11916;
  wire       [15:0]   _zz_11917;
  wire       [15:0]   _zz_11918;
  wire       [15:0]   _zz_11919;
  wire       [15:0]   _zz_11920;
  wire       [15:0]   _zz_11921;
  wire       [15:0]   _zz_11922;
  wire       [15:0]   _zz_11923;
  wire       [15:0]   _zz_11924;
  wire       [15:0]   _zz_11925;
  wire       [15:0]   _zz_11926;
  wire       [15:0]   _zz_11927;
  wire       [15:0]   _zz_11928;
  wire       [15:0]   _zz_11929;
  wire       [15:0]   _zz_11930;
  wire       [31:0]   _zz_11931;
  wire       [31:0]   _zz_11932;
  wire       [15:0]   _zz_11933;
  wire       [31:0]   _zz_11934;
  wire       [31:0]   _zz_11935;
  wire       [15:0]   _zz_11936;
  wire       [15:0]   _zz_11937;
  wire       [15:0]   _zz_11938;
  wire       [15:0]   _zz_11939;
  wire       [15:0]   _zz_11940;
  wire       [15:0]   _zz_11941;
  wire       [15:0]   _zz_11942;
  wire       [15:0]   _zz_11943;
  wire       [15:0]   _zz_11944;
  wire       [15:0]   _zz_11945;
  wire       [15:0]   _zz_11946;
  wire       [15:0]   _zz_11947;
  wire       [15:0]   _zz_11948;
  wire       [15:0]   _zz_11949;
  wire       [15:0]   _zz_11950;
  wire       [15:0]   _zz_11951;
  wire       [15:0]   _zz_11952;
  wire       [31:0]   _zz_11953;
  wire       [31:0]   _zz_11954;
  wire       [15:0]   _zz_11955;
  wire       [31:0]   _zz_11956;
  wire       [31:0]   _zz_11957;
  wire       [15:0]   _zz_11958;
  wire       [15:0]   _zz_11959;
  wire       [15:0]   _zz_11960;
  wire       [15:0]   _zz_11961;
  wire       [15:0]   _zz_11962;
  wire       [15:0]   _zz_11963;
  wire       [15:0]   _zz_11964;
  wire       [15:0]   _zz_11965;
  wire       [15:0]   _zz_11966;
  wire       [15:0]   _zz_11967;
  wire       [15:0]   _zz_11968;
  wire       [15:0]   _zz_11969;
  wire       [15:0]   _zz_11970;
  wire       [15:0]   _zz_11971;
  wire       [15:0]   _zz_11972;
  wire       [15:0]   _zz_11973;
  wire       [15:0]   _zz_11974;
  wire       [31:0]   _zz_11975;
  wire       [31:0]   _zz_11976;
  wire       [15:0]   _zz_11977;
  wire       [31:0]   _zz_11978;
  wire       [31:0]   _zz_11979;
  wire       [15:0]   _zz_11980;
  wire       [15:0]   _zz_11981;
  wire       [15:0]   _zz_11982;
  wire       [15:0]   _zz_11983;
  wire       [15:0]   _zz_11984;
  wire       [15:0]   _zz_11985;
  wire       [15:0]   _zz_11986;
  wire       [15:0]   _zz_11987;
  wire       [15:0]   _zz_11988;
  wire       [15:0]   _zz_11989;
  wire       [15:0]   _zz_11990;
  wire       [15:0]   _zz_11991;
  wire       [15:0]   _zz_11992;
  wire       [15:0]   _zz_11993;
  wire       [15:0]   _zz_11994;
  wire       [15:0]   _zz_11995;
  wire       [15:0]   _zz_11996;
  wire       [31:0]   _zz_11997;
  wire       [31:0]   _zz_11998;
  wire       [15:0]   _zz_11999;
  wire       [31:0]   _zz_12000;
  wire       [31:0]   _zz_12001;
  wire       [15:0]   _zz_12002;
  wire       [15:0]   _zz_12003;
  wire       [15:0]   _zz_12004;
  wire       [15:0]   _zz_12005;
  wire       [15:0]   _zz_12006;
  wire       [15:0]   _zz_12007;
  wire       [15:0]   _zz_12008;
  wire       [15:0]   _zz_12009;
  wire       [15:0]   _zz_12010;
  wire       [15:0]   _zz_12011;
  wire       [15:0]   _zz_12012;
  wire       [15:0]   _zz_12013;
  wire       [15:0]   _zz_12014;
  wire       [15:0]   _zz_12015;
  wire       [15:0]   _zz_12016;
  wire       [15:0]   _zz_12017;
  wire       [15:0]   _zz_12018;
  wire       [31:0]   _zz_12019;
  wire       [31:0]   _zz_12020;
  wire       [15:0]   _zz_12021;
  wire       [31:0]   _zz_12022;
  wire       [31:0]   _zz_12023;
  wire       [15:0]   _zz_12024;
  wire       [15:0]   _zz_12025;
  wire       [15:0]   _zz_12026;
  wire       [15:0]   _zz_12027;
  wire       [15:0]   _zz_12028;
  wire       [15:0]   _zz_12029;
  wire       [15:0]   _zz_12030;
  wire       [15:0]   _zz_12031;
  wire       [15:0]   _zz_12032;
  wire       [15:0]   _zz_12033;
  wire       [15:0]   _zz_12034;
  wire       [15:0]   _zz_12035;
  wire       [15:0]   _zz_12036;
  wire       [15:0]   _zz_12037;
  wire       [15:0]   _zz_12038;
  wire       [15:0]   _zz_12039;
  wire       [15:0]   _zz_12040;
  wire       [31:0]   _zz_12041;
  wire       [31:0]   _zz_12042;
  wire       [15:0]   _zz_12043;
  wire       [31:0]   _zz_12044;
  wire       [31:0]   _zz_12045;
  wire       [15:0]   _zz_12046;
  wire       [15:0]   _zz_12047;
  wire       [15:0]   _zz_12048;
  wire       [15:0]   _zz_12049;
  wire       [15:0]   _zz_12050;
  wire       [15:0]   _zz_12051;
  wire       [15:0]   _zz_12052;
  wire       [15:0]   _zz_12053;
  wire       [15:0]   _zz_12054;
  wire       [15:0]   _zz_12055;
  wire       [15:0]   _zz_12056;
  wire       [15:0]   _zz_12057;
  wire       [15:0]   _zz_12058;
  wire       [15:0]   _zz_12059;
  wire       [15:0]   _zz_12060;
  wire       [15:0]   _zz_12061;
  wire       [15:0]   _zz_12062;
  wire       [31:0]   _zz_12063;
  wire       [31:0]   _zz_12064;
  wire       [15:0]   _zz_12065;
  wire       [31:0]   _zz_12066;
  wire       [31:0]   _zz_12067;
  wire       [15:0]   _zz_12068;
  wire       [15:0]   _zz_12069;
  wire       [15:0]   _zz_12070;
  wire       [15:0]   _zz_12071;
  wire       [15:0]   _zz_12072;
  wire       [15:0]   _zz_12073;
  wire       [15:0]   _zz_12074;
  wire       [15:0]   _zz_12075;
  wire       [15:0]   _zz_12076;
  wire       [15:0]   _zz_12077;
  wire       [15:0]   _zz_12078;
  wire       [15:0]   _zz_12079;
  wire       [15:0]   _zz_12080;
  wire       [15:0]   _zz_12081;
  wire       [15:0]   _zz_12082;
  wire       [15:0]   _zz_12083;
  wire       [15:0]   _zz_12084;
  wire       [31:0]   _zz_12085;
  wire       [31:0]   _zz_12086;
  wire       [15:0]   _zz_12087;
  wire       [31:0]   _zz_12088;
  wire       [31:0]   _zz_12089;
  wire       [15:0]   _zz_12090;
  wire       [15:0]   _zz_12091;
  wire       [15:0]   _zz_12092;
  wire       [15:0]   _zz_12093;
  wire       [15:0]   _zz_12094;
  wire       [15:0]   _zz_12095;
  wire       [15:0]   _zz_12096;
  wire       [15:0]   _zz_12097;
  wire       [15:0]   _zz_12098;
  wire       [15:0]   _zz_12099;
  wire       [15:0]   _zz_12100;
  wire       [15:0]   _zz_12101;
  wire       [15:0]   _zz_12102;
  wire       [15:0]   _zz_12103;
  wire       [15:0]   _zz_12104;
  wire       [15:0]   _zz_12105;
  wire       [15:0]   _zz_12106;
  wire       [31:0]   _zz_12107;
  wire       [31:0]   _zz_12108;
  wire       [15:0]   _zz_12109;
  wire       [31:0]   _zz_12110;
  wire       [31:0]   _zz_12111;
  wire       [15:0]   _zz_12112;
  wire       [15:0]   _zz_12113;
  wire       [15:0]   _zz_12114;
  wire       [15:0]   _zz_12115;
  wire       [15:0]   _zz_12116;
  wire       [15:0]   _zz_12117;
  wire       [15:0]   _zz_12118;
  wire       [15:0]   _zz_12119;
  wire       [15:0]   _zz_12120;
  wire       [15:0]   _zz_12121;
  wire       [15:0]   _zz_12122;
  wire       [15:0]   _zz_12123;
  wire       [15:0]   _zz_12124;
  wire       [15:0]   _zz_12125;
  wire       [15:0]   _zz_12126;
  wire       [15:0]   _zz_12127;
  wire       [15:0]   _zz_12128;
  wire       [31:0]   _zz_12129;
  wire       [31:0]   _zz_12130;
  wire       [15:0]   _zz_12131;
  wire       [31:0]   _zz_12132;
  wire       [31:0]   _zz_12133;
  wire       [15:0]   _zz_12134;
  wire       [15:0]   _zz_12135;
  wire       [15:0]   _zz_12136;
  wire       [15:0]   _zz_12137;
  wire       [15:0]   _zz_12138;
  wire       [15:0]   _zz_12139;
  wire       [15:0]   _zz_12140;
  wire       [15:0]   _zz_12141;
  wire       [15:0]   _zz_12142;
  wire       [15:0]   _zz_12143;
  wire       [15:0]   _zz_12144;
  wire       [15:0]   _zz_12145;
  wire       [15:0]   _zz_12146;
  wire       [15:0]   _zz_12147;
  wire       [15:0]   _zz_12148;
  wire       [15:0]   _zz_12149;
  wire       [15:0]   _zz_12150;
  wire       [31:0]   _zz_12151;
  wire       [31:0]   _zz_12152;
  wire       [15:0]   _zz_12153;
  wire       [31:0]   _zz_12154;
  wire       [31:0]   _zz_12155;
  wire       [15:0]   _zz_12156;
  wire       [15:0]   _zz_12157;
  wire       [15:0]   _zz_12158;
  wire       [15:0]   _zz_12159;
  wire       [15:0]   _zz_12160;
  wire       [15:0]   _zz_12161;
  wire       [15:0]   _zz_12162;
  wire       [15:0]   _zz_12163;
  wire       [15:0]   _zz_12164;
  wire       [15:0]   _zz_12165;
  wire       [15:0]   _zz_12166;
  wire       [15:0]   _zz_12167;
  wire       [15:0]   _zz_12168;
  wire       [15:0]   _zz_12169;
  wire       [15:0]   _zz_12170;
  wire       [15:0]   _zz_12171;
  wire       [15:0]   _zz_12172;
  wire       [31:0]   _zz_12173;
  wire       [31:0]   _zz_12174;
  wire       [15:0]   _zz_12175;
  wire       [31:0]   _zz_12176;
  wire       [31:0]   _zz_12177;
  wire       [15:0]   _zz_12178;
  wire       [15:0]   _zz_12179;
  wire       [15:0]   _zz_12180;
  wire       [15:0]   _zz_12181;
  wire       [15:0]   _zz_12182;
  wire       [15:0]   _zz_12183;
  wire       [15:0]   _zz_12184;
  wire       [15:0]   _zz_12185;
  wire       [15:0]   _zz_12186;
  wire       [15:0]   _zz_12187;
  wire       [15:0]   _zz_12188;
  wire       [15:0]   _zz_12189;
  wire       [15:0]   _zz_12190;
  wire       [15:0]   _zz_12191;
  wire       [15:0]   _zz_12192;
  wire       [15:0]   _zz_12193;
  wire       [15:0]   _zz_12194;
  wire       [31:0]   _zz_12195;
  wire       [31:0]   _zz_12196;
  wire       [15:0]   _zz_12197;
  wire       [31:0]   _zz_12198;
  wire       [31:0]   _zz_12199;
  wire       [15:0]   _zz_12200;
  wire       [15:0]   _zz_12201;
  wire       [15:0]   _zz_12202;
  wire       [15:0]   _zz_12203;
  wire       [15:0]   _zz_12204;
  wire       [15:0]   _zz_12205;
  wire       [15:0]   _zz_12206;
  wire       [15:0]   _zz_12207;
  wire       [15:0]   _zz_12208;
  wire       [15:0]   _zz_12209;
  wire       [15:0]   _zz_12210;
  wire       [15:0]   _zz_12211;
  wire       [15:0]   _zz_12212;
  wire       [15:0]   _zz_12213;
  wire       [15:0]   _zz_12214;
  wire       [15:0]   _zz_12215;
  wire       [15:0]   _zz_12216;
  wire       [31:0]   _zz_12217;
  wire       [31:0]   _zz_12218;
  wire       [15:0]   _zz_12219;
  wire       [31:0]   _zz_12220;
  wire       [31:0]   _zz_12221;
  wire       [15:0]   _zz_12222;
  wire       [15:0]   _zz_12223;
  wire       [15:0]   _zz_12224;
  wire       [15:0]   _zz_12225;
  wire       [15:0]   _zz_12226;
  wire       [15:0]   _zz_12227;
  wire       [15:0]   _zz_12228;
  wire       [15:0]   _zz_12229;
  wire       [15:0]   _zz_12230;
  wire       [15:0]   _zz_12231;
  wire       [15:0]   _zz_12232;
  wire       [15:0]   _zz_12233;
  wire       [15:0]   _zz_12234;
  wire       [15:0]   _zz_12235;
  wire       [15:0]   _zz_12236;
  wire       [15:0]   _zz_12237;
  wire       [15:0]   _zz_12238;
  wire       [31:0]   _zz_12239;
  wire       [31:0]   _zz_12240;
  wire       [15:0]   _zz_12241;
  wire       [31:0]   _zz_12242;
  wire       [31:0]   _zz_12243;
  wire       [15:0]   _zz_12244;
  wire       [15:0]   _zz_12245;
  wire       [15:0]   _zz_12246;
  wire       [15:0]   _zz_12247;
  wire       [15:0]   _zz_12248;
  wire       [15:0]   _zz_12249;
  wire       [15:0]   _zz_12250;
  wire       [15:0]   _zz_12251;
  wire       [15:0]   _zz_12252;
  wire       [15:0]   _zz_12253;
  wire       [15:0]   _zz_12254;
  wire       [15:0]   _zz_12255;
  wire       [15:0]   _zz_12256;
  wire       [15:0]   _zz_12257;
  wire       [15:0]   _zz_12258;
  wire       [15:0]   _zz_12259;
  wire       [15:0]   _zz_12260;
  wire       [31:0]   _zz_12261;
  wire       [31:0]   _zz_12262;
  wire       [15:0]   _zz_12263;
  wire       [31:0]   _zz_12264;
  wire       [31:0]   _zz_12265;
  wire       [15:0]   _zz_12266;
  wire       [15:0]   _zz_12267;
  wire       [15:0]   _zz_12268;
  wire       [15:0]   _zz_12269;
  wire       [15:0]   _zz_12270;
  wire       [15:0]   _zz_12271;
  wire       [15:0]   _zz_12272;
  wire       [15:0]   _zz_12273;
  wire       [15:0]   _zz_12274;
  wire       [15:0]   _zz_12275;
  wire       [15:0]   _zz_12276;
  wire       [15:0]   _zz_12277;
  wire       [15:0]   _zz_12278;
  wire       [15:0]   _zz_12279;
  wire       [15:0]   _zz_12280;
  wire       [15:0]   _zz_12281;
  wire       [15:0]   _zz_12282;
  wire       [31:0]   _zz_12283;
  wire       [31:0]   _zz_12284;
  wire       [15:0]   _zz_12285;
  wire       [31:0]   _zz_12286;
  wire       [31:0]   _zz_12287;
  wire       [15:0]   _zz_12288;
  wire       [15:0]   _zz_12289;
  wire       [15:0]   _zz_12290;
  wire       [15:0]   _zz_12291;
  wire       [15:0]   _zz_12292;
  wire       [15:0]   _zz_12293;
  wire       [15:0]   _zz_12294;
  wire       [15:0]   _zz_12295;
  wire       [15:0]   _zz_12296;
  wire       [15:0]   _zz_12297;
  wire       [15:0]   _zz_12298;
  wire       [15:0]   _zz_12299;
  wire       [15:0]   _zz_12300;
  wire       [15:0]   _zz_12301;
  wire       [15:0]   _zz_12302;
  wire       [15:0]   _zz_12303;
  wire       [15:0]   _zz_12304;
  wire       [31:0]   _zz_12305;
  wire       [31:0]   _zz_12306;
  wire       [15:0]   _zz_12307;
  wire       [31:0]   _zz_12308;
  wire       [31:0]   _zz_12309;
  wire       [15:0]   _zz_12310;
  wire       [15:0]   _zz_12311;
  wire       [15:0]   _zz_12312;
  wire       [15:0]   _zz_12313;
  wire       [15:0]   _zz_12314;
  wire       [15:0]   _zz_12315;
  wire       [15:0]   _zz_12316;
  wire       [15:0]   _zz_12317;
  wire       [15:0]   _zz_12318;
  wire       [15:0]   _zz_12319;
  wire       [15:0]   _zz_12320;
  wire       [15:0]   _zz_12321;
  wire       [15:0]   _zz_12322;
  wire       [15:0]   _zz_12323;
  wire       [15:0]   _zz_12324;
  wire       [15:0]   _zz_12325;
  wire       [15:0]   _zz_12326;
  wire       [31:0]   _zz_12327;
  wire       [31:0]   _zz_12328;
  wire       [15:0]   _zz_12329;
  wire       [31:0]   _zz_12330;
  wire       [31:0]   _zz_12331;
  wire       [15:0]   _zz_12332;
  wire       [15:0]   _zz_12333;
  wire       [15:0]   _zz_12334;
  wire       [15:0]   _zz_12335;
  wire       [15:0]   _zz_12336;
  wire       [15:0]   _zz_12337;
  wire       [15:0]   _zz_12338;
  wire       [15:0]   _zz_12339;
  wire       [15:0]   _zz_12340;
  wire       [15:0]   _zz_12341;
  wire       [15:0]   _zz_12342;
  wire       [15:0]   _zz_12343;
  wire       [15:0]   _zz_12344;
  wire       [15:0]   _zz_12345;
  wire       [15:0]   _zz_12346;
  wire       [15:0]   _zz_12347;
  wire       [15:0]   _zz_12348;
  wire       [31:0]   _zz_12349;
  wire       [31:0]   _zz_12350;
  wire       [15:0]   _zz_12351;
  wire       [31:0]   _zz_12352;
  wire       [31:0]   _zz_12353;
  wire       [15:0]   _zz_12354;
  wire       [15:0]   _zz_12355;
  wire       [15:0]   _zz_12356;
  wire       [15:0]   _zz_12357;
  wire       [15:0]   _zz_12358;
  wire       [15:0]   _zz_12359;
  wire       [15:0]   _zz_12360;
  wire       [15:0]   _zz_12361;
  wire       [15:0]   _zz_12362;
  wire       [15:0]   _zz_12363;
  wire       [15:0]   _zz_12364;
  wire       [15:0]   _zz_12365;
  wire       [15:0]   _zz_12366;
  wire       [15:0]   _zz_12367;
  wire       [15:0]   _zz_12368;
  wire       [15:0]   _zz_12369;
  wire       [15:0]   _zz_12370;
  wire       [31:0]   _zz_12371;
  wire       [31:0]   _zz_12372;
  wire       [15:0]   _zz_12373;
  wire       [31:0]   _zz_12374;
  wire       [31:0]   _zz_12375;
  wire       [15:0]   _zz_12376;
  wire       [15:0]   _zz_12377;
  wire       [15:0]   _zz_12378;
  wire       [15:0]   _zz_12379;
  wire       [15:0]   _zz_12380;
  wire       [15:0]   _zz_12381;
  wire       [15:0]   _zz_12382;
  wire       [15:0]   _zz_12383;
  wire       [15:0]   _zz_12384;
  wire       [15:0]   _zz_12385;
  wire       [15:0]   _zz_12386;
  wire       [15:0]   _zz_12387;
  wire       [15:0]   _zz_12388;
  wire       [15:0]   _zz_12389;
  wire       [15:0]   _zz_12390;
  wire       [15:0]   _zz_12391;
  wire       [15:0]   _zz_12392;
  wire       [31:0]   _zz_12393;
  wire       [31:0]   _zz_12394;
  wire       [15:0]   _zz_12395;
  wire       [31:0]   _zz_12396;
  wire       [31:0]   _zz_12397;
  wire       [15:0]   _zz_12398;
  wire       [15:0]   _zz_12399;
  wire       [15:0]   _zz_12400;
  wire       [15:0]   _zz_12401;
  wire       [15:0]   _zz_12402;
  wire       [15:0]   _zz_12403;
  wire       [15:0]   _zz_12404;
  wire       [15:0]   _zz_12405;
  wire       [15:0]   _zz_12406;
  wire       [15:0]   _zz_12407;
  wire       [15:0]   _zz_12408;
  wire       [15:0]   _zz_12409;
  wire       [15:0]   _zz_12410;
  wire       [15:0]   _zz_12411;
  wire       [15:0]   _zz_12412;
  wire       [15:0]   _zz_12413;
  wire       [15:0]   _zz_12414;
  wire       [31:0]   _zz_12415;
  wire       [31:0]   _zz_12416;
  wire       [15:0]   _zz_12417;
  wire       [31:0]   _zz_12418;
  wire       [31:0]   _zz_12419;
  wire       [15:0]   _zz_12420;
  wire       [15:0]   _zz_12421;
  wire       [15:0]   _zz_12422;
  wire       [15:0]   _zz_12423;
  wire       [15:0]   _zz_12424;
  wire       [15:0]   _zz_12425;
  wire       [15:0]   _zz_12426;
  wire       [15:0]   _zz_12427;
  wire       [15:0]   _zz_12428;
  wire       [15:0]   _zz_12429;
  wire       [15:0]   _zz_12430;
  wire       [15:0]   _zz_12431;
  wire       [15:0]   _zz_12432;
  wire       [15:0]   _zz_12433;
  wire       [15:0]   _zz_12434;
  wire       [15:0]   _zz_12435;
  wire       [15:0]   _zz_12436;
  wire       [31:0]   _zz_12437;
  wire       [31:0]   _zz_12438;
  wire       [15:0]   _zz_12439;
  wire       [31:0]   _zz_12440;
  wire       [31:0]   _zz_12441;
  wire       [15:0]   _zz_12442;
  wire       [15:0]   _zz_12443;
  wire       [15:0]   _zz_12444;
  wire       [15:0]   _zz_12445;
  wire       [15:0]   _zz_12446;
  wire       [15:0]   _zz_12447;
  wire       [15:0]   _zz_12448;
  wire       [15:0]   _zz_12449;
  wire       [15:0]   _zz_12450;
  wire       [15:0]   _zz_12451;
  wire       [15:0]   _zz_12452;
  wire       [15:0]   _zz_12453;
  wire       [15:0]   _zz_12454;
  wire       [15:0]   _zz_12455;
  wire       [15:0]   _zz_12456;
  wire       [15:0]   _zz_12457;
  wire       [15:0]   _zz_12458;
  wire       [31:0]   _zz_12459;
  wire       [31:0]   _zz_12460;
  wire       [15:0]   _zz_12461;
  wire       [31:0]   _zz_12462;
  wire       [31:0]   _zz_12463;
  wire       [15:0]   _zz_12464;
  wire       [15:0]   _zz_12465;
  wire       [15:0]   _zz_12466;
  wire       [15:0]   _zz_12467;
  wire       [15:0]   _zz_12468;
  wire       [15:0]   _zz_12469;
  wire       [15:0]   _zz_12470;
  wire       [15:0]   _zz_12471;
  wire       [15:0]   _zz_12472;
  wire       [15:0]   _zz_12473;
  wire       [15:0]   _zz_12474;
  wire       [15:0]   _zz_12475;
  wire       [15:0]   _zz_12476;
  wire       [15:0]   _zz_12477;
  wire       [15:0]   _zz_12478;
  wire       [15:0]   _zz_12479;
  wire       [15:0]   _zz_12480;
  wire       [31:0]   _zz_12481;
  wire       [31:0]   _zz_12482;
  wire       [15:0]   _zz_12483;
  wire       [31:0]   _zz_12484;
  wire       [31:0]   _zz_12485;
  wire       [15:0]   _zz_12486;
  wire       [15:0]   _zz_12487;
  wire       [15:0]   _zz_12488;
  wire       [15:0]   _zz_12489;
  wire       [15:0]   _zz_12490;
  wire       [15:0]   _zz_12491;
  wire       [15:0]   _zz_12492;
  wire       [15:0]   _zz_12493;
  wire       [15:0]   _zz_12494;
  wire       [15:0]   _zz_12495;
  wire       [15:0]   _zz_12496;
  wire       [15:0]   _zz_12497;
  wire       [15:0]   _zz_12498;
  wire       [15:0]   _zz_12499;
  wire       [15:0]   _zz_12500;
  wire       [15:0]   _zz_12501;
  wire       [15:0]   _zz_12502;
  wire       [31:0]   _zz_12503;
  wire       [31:0]   _zz_12504;
  wire       [15:0]   _zz_12505;
  wire       [31:0]   _zz_12506;
  wire       [31:0]   _zz_12507;
  wire       [15:0]   _zz_12508;
  wire       [15:0]   _zz_12509;
  wire       [15:0]   _zz_12510;
  wire       [15:0]   _zz_12511;
  wire       [15:0]   _zz_12512;
  wire       [15:0]   _zz_12513;
  wire       [15:0]   _zz_12514;
  wire       [15:0]   _zz_12515;
  wire       [15:0]   _zz_12516;
  wire       [15:0]   _zz_12517;
  wire       [15:0]   _zz_12518;
  wire       [15:0]   _zz_12519;
  wire       [15:0]   _zz_12520;
  wire       [15:0]   _zz_12521;
  wire       [15:0]   _zz_12522;
  wire       [15:0]   _zz_12523;
  wire       [15:0]   _zz_12524;
  wire       [31:0]   _zz_12525;
  wire       [31:0]   _zz_12526;
  wire       [15:0]   _zz_12527;
  wire       [31:0]   _zz_12528;
  wire       [31:0]   _zz_12529;
  wire       [15:0]   _zz_12530;
  wire       [15:0]   _zz_12531;
  wire       [15:0]   _zz_12532;
  wire       [15:0]   _zz_12533;
  wire       [15:0]   _zz_12534;
  wire       [15:0]   _zz_12535;
  wire       [15:0]   _zz_12536;
  wire       [15:0]   _zz_12537;
  wire       [15:0]   _zz_12538;
  wire       [15:0]   _zz_12539;
  wire       [15:0]   _zz_12540;
  wire       [15:0]   _zz_12541;
  wire       [15:0]   _zz_12542;
  wire       [15:0]   _zz_12543;
  wire       [15:0]   _zz_12544;
  wire       [15:0]   _zz_12545;
  wire       [15:0]   _zz_12546;
  reg        [15:0]   data_in_0_real;
  reg        [15:0]   data_in_0_imag;
  reg        [15:0]   data_in_1_real;
  reg        [15:0]   data_in_1_imag;
  reg        [15:0]   data_in_2_real;
  reg        [15:0]   data_in_2_imag;
  reg        [15:0]   data_in_3_real;
  reg        [15:0]   data_in_3_imag;
  reg        [15:0]   data_in_4_real;
  reg        [15:0]   data_in_4_imag;
  reg        [15:0]   data_in_5_real;
  reg        [15:0]   data_in_5_imag;
  reg        [15:0]   data_in_6_real;
  reg        [15:0]   data_in_6_imag;
  reg        [15:0]   data_in_7_real;
  reg        [15:0]   data_in_7_imag;
  reg        [15:0]   data_in_8_real;
  reg        [15:0]   data_in_8_imag;
  reg        [15:0]   data_in_9_real;
  reg        [15:0]   data_in_9_imag;
  reg        [15:0]   data_in_10_real;
  reg        [15:0]   data_in_10_imag;
  reg        [15:0]   data_in_11_real;
  reg        [15:0]   data_in_11_imag;
  reg        [15:0]   data_in_12_real;
  reg        [15:0]   data_in_12_imag;
  reg        [15:0]   data_in_13_real;
  reg        [15:0]   data_in_13_imag;
  reg        [15:0]   data_in_14_real;
  reg        [15:0]   data_in_14_imag;
  reg        [15:0]   data_in_15_real;
  reg        [15:0]   data_in_15_imag;
  reg        [15:0]   data_in_16_real;
  reg        [15:0]   data_in_16_imag;
  reg        [15:0]   data_in_17_real;
  reg        [15:0]   data_in_17_imag;
  reg        [15:0]   data_in_18_real;
  reg        [15:0]   data_in_18_imag;
  reg        [15:0]   data_in_19_real;
  reg        [15:0]   data_in_19_imag;
  reg        [15:0]   data_in_20_real;
  reg        [15:0]   data_in_20_imag;
  reg        [15:0]   data_in_21_real;
  reg        [15:0]   data_in_21_imag;
  reg        [15:0]   data_in_22_real;
  reg        [15:0]   data_in_22_imag;
  reg        [15:0]   data_in_23_real;
  reg        [15:0]   data_in_23_imag;
  reg        [15:0]   data_in_24_real;
  reg        [15:0]   data_in_24_imag;
  reg        [15:0]   data_in_25_real;
  reg        [15:0]   data_in_25_imag;
  reg        [15:0]   data_in_26_real;
  reg        [15:0]   data_in_26_imag;
  reg        [15:0]   data_in_27_real;
  reg        [15:0]   data_in_27_imag;
  reg        [15:0]   data_in_28_real;
  reg        [15:0]   data_in_28_imag;
  reg        [15:0]   data_in_29_real;
  reg        [15:0]   data_in_29_imag;
  reg        [15:0]   data_in_30_real;
  reg        [15:0]   data_in_30_imag;
  reg        [15:0]   data_in_31_real;
  reg        [15:0]   data_in_31_imag;
  reg        [15:0]   data_in_32_real;
  reg        [15:0]   data_in_32_imag;
  reg        [15:0]   data_in_33_real;
  reg        [15:0]   data_in_33_imag;
  reg        [15:0]   data_in_34_real;
  reg        [15:0]   data_in_34_imag;
  reg        [15:0]   data_in_35_real;
  reg        [15:0]   data_in_35_imag;
  reg        [15:0]   data_in_36_real;
  reg        [15:0]   data_in_36_imag;
  reg        [15:0]   data_in_37_real;
  reg        [15:0]   data_in_37_imag;
  reg        [15:0]   data_in_38_real;
  reg        [15:0]   data_in_38_imag;
  reg        [15:0]   data_in_39_real;
  reg        [15:0]   data_in_39_imag;
  reg        [15:0]   data_in_40_real;
  reg        [15:0]   data_in_40_imag;
  reg        [15:0]   data_in_41_real;
  reg        [15:0]   data_in_41_imag;
  reg        [15:0]   data_in_42_real;
  reg        [15:0]   data_in_42_imag;
  reg        [15:0]   data_in_43_real;
  reg        [15:0]   data_in_43_imag;
  reg        [15:0]   data_in_44_real;
  reg        [15:0]   data_in_44_imag;
  reg        [15:0]   data_in_45_real;
  reg        [15:0]   data_in_45_imag;
  reg        [15:0]   data_in_46_real;
  reg        [15:0]   data_in_46_imag;
  reg        [15:0]   data_in_47_real;
  reg        [15:0]   data_in_47_imag;
  reg        [15:0]   data_in_48_real;
  reg        [15:0]   data_in_48_imag;
  reg        [15:0]   data_in_49_real;
  reg        [15:0]   data_in_49_imag;
  reg        [15:0]   data_in_50_real;
  reg        [15:0]   data_in_50_imag;
  reg        [15:0]   data_in_51_real;
  reg        [15:0]   data_in_51_imag;
  reg        [15:0]   data_in_52_real;
  reg        [15:0]   data_in_52_imag;
  reg        [15:0]   data_in_53_real;
  reg        [15:0]   data_in_53_imag;
  reg        [15:0]   data_in_54_real;
  reg        [15:0]   data_in_54_imag;
  reg        [15:0]   data_in_55_real;
  reg        [15:0]   data_in_55_imag;
  reg        [15:0]   data_in_56_real;
  reg        [15:0]   data_in_56_imag;
  reg        [15:0]   data_in_57_real;
  reg        [15:0]   data_in_57_imag;
  reg        [15:0]   data_in_58_real;
  reg        [15:0]   data_in_58_imag;
  reg        [15:0]   data_in_59_real;
  reg        [15:0]   data_in_59_imag;
  reg        [15:0]   data_in_60_real;
  reg        [15:0]   data_in_60_imag;
  reg        [15:0]   data_in_61_real;
  reg        [15:0]   data_in_61_imag;
  reg        [15:0]   data_in_62_real;
  reg        [15:0]   data_in_62_imag;
  reg        [15:0]   data_in_63_real;
  reg        [15:0]   data_in_63_imag;
  reg        [15:0]   data_in_64_real;
  reg        [15:0]   data_in_64_imag;
  reg        [15:0]   data_in_65_real;
  reg        [15:0]   data_in_65_imag;
  reg        [15:0]   data_in_66_real;
  reg        [15:0]   data_in_66_imag;
  reg        [15:0]   data_in_67_real;
  reg        [15:0]   data_in_67_imag;
  reg        [15:0]   data_in_68_real;
  reg        [15:0]   data_in_68_imag;
  reg        [15:0]   data_in_69_real;
  reg        [15:0]   data_in_69_imag;
  reg        [15:0]   data_in_70_real;
  reg        [15:0]   data_in_70_imag;
  reg        [15:0]   data_in_71_real;
  reg        [15:0]   data_in_71_imag;
  reg        [15:0]   data_in_72_real;
  reg        [15:0]   data_in_72_imag;
  reg        [15:0]   data_in_73_real;
  reg        [15:0]   data_in_73_imag;
  reg        [15:0]   data_in_74_real;
  reg        [15:0]   data_in_74_imag;
  reg        [15:0]   data_in_75_real;
  reg        [15:0]   data_in_75_imag;
  reg        [15:0]   data_in_76_real;
  reg        [15:0]   data_in_76_imag;
  reg        [15:0]   data_in_77_real;
  reg        [15:0]   data_in_77_imag;
  reg        [15:0]   data_in_78_real;
  reg        [15:0]   data_in_78_imag;
  reg        [15:0]   data_in_79_real;
  reg        [15:0]   data_in_79_imag;
  reg        [15:0]   data_in_80_real;
  reg        [15:0]   data_in_80_imag;
  reg        [15:0]   data_in_81_real;
  reg        [15:0]   data_in_81_imag;
  reg        [15:0]   data_in_82_real;
  reg        [15:0]   data_in_82_imag;
  reg        [15:0]   data_in_83_real;
  reg        [15:0]   data_in_83_imag;
  reg        [15:0]   data_in_84_real;
  reg        [15:0]   data_in_84_imag;
  reg        [15:0]   data_in_85_real;
  reg        [15:0]   data_in_85_imag;
  reg        [15:0]   data_in_86_real;
  reg        [15:0]   data_in_86_imag;
  reg        [15:0]   data_in_87_real;
  reg        [15:0]   data_in_87_imag;
  reg        [15:0]   data_in_88_real;
  reg        [15:0]   data_in_88_imag;
  reg        [15:0]   data_in_89_real;
  reg        [15:0]   data_in_89_imag;
  reg        [15:0]   data_in_90_real;
  reg        [15:0]   data_in_90_imag;
  reg        [15:0]   data_in_91_real;
  reg        [15:0]   data_in_91_imag;
  reg        [15:0]   data_in_92_real;
  reg        [15:0]   data_in_92_imag;
  reg        [15:0]   data_in_93_real;
  reg        [15:0]   data_in_93_imag;
  reg        [15:0]   data_in_94_real;
  reg        [15:0]   data_in_94_imag;
  reg        [15:0]   data_in_95_real;
  reg        [15:0]   data_in_95_imag;
  reg        [15:0]   data_in_96_real;
  reg        [15:0]   data_in_96_imag;
  reg        [15:0]   data_in_97_real;
  reg        [15:0]   data_in_97_imag;
  reg        [15:0]   data_in_98_real;
  reg        [15:0]   data_in_98_imag;
  reg        [15:0]   data_in_99_real;
  reg        [15:0]   data_in_99_imag;
  reg        [15:0]   data_in_100_real;
  reg        [15:0]   data_in_100_imag;
  reg        [15:0]   data_in_101_real;
  reg        [15:0]   data_in_101_imag;
  reg        [15:0]   data_in_102_real;
  reg        [15:0]   data_in_102_imag;
  reg        [15:0]   data_in_103_real;
  reg        [15:0]   data_in_103_imag;
  reg        [15:0]   data_in_104_real;
  reg        [15:0]   data_in_104_imag;
  reg        [15:0]   data_in_105_real;
  reg        [15:0]   data_in_105_imag;
  reg        [15:0]   data_in_106_real;
  reg        [15:0]   data_in_106_imag;
  reg        [15:0]   data_in_107_real;
  reg        [15:0]   data_in_107_imag;
  reg        [15:0]   data_in_108_real;
  reg        [15:0]   data_in_108_imag;
  reg        [15:0]   data_in_109_real;
  reg        [15:0]   data_in_109_imag;
  reg        [15:0]   data_in_110_real;
  reg        [15:0]   data_in_110_imag;
  reg        [15:0]   data_in_111_real;
  reg        [15:0]   data_in_111_imag;
  reg        [15:0]   data_in_112_real;
  reg        [15:0]   data_in_112_imag;
  reg        [15:0]   data_in_113_real;
  reg        [15:0]   data_in_113_imag;
  reg        [15:0]   data_in_114_real;
  reg        [15:0]   data_in_114_imag;
  reg        [15:0]   data_in_115_real;
  reg        [15:0]   data_in_115_imag;
  reg        [15:0]   data_in_116_real;
  reg        [15:0]   data_in_116_imag;
  reg        [15:0]   data_in_117_real;
  reg        [15:0]   data_in_117_imag;
  reg        [15:0]   data_in_118_real;
  reg        [15:0]   data_in_118_imag;
  reg        [15:0]   data_in_119_real;
  reg        [15:0]   data_in_119_imag;
  reg        [15:0]   data_in_120_real;
  reg        [15:0]   data_in_120_imag;
  reg        [15:0]   data_in_121_real;
  reg        [15:0]   data_in_121_imag;
  reg        [15:0]   data_in_122_real;
  reg        [15:0]   data_in_122_imag;
  reg        [15:0]   data_in_123_real;
  reg        [15:0]   data_in_123_imag;
  reg        [15:0]   data_in_124_real;
  reg        [15:0]   data_in_124_imag;
  reg        [15:0]   data_in_125_real;
  reg        [15:0]   data_in_125_imag;
  reg        [15:0]   data_in_126_real;
  reg        [15:0]   data_in_126_imag;
  reg        [15:0]   data_in_127_real;
  reg        [15:0]   data_in_127_imag;
  wire       [15:0]   twiddle_factor_table_0_real;
  wire       [15:0]   twiddle_factor_table_0_imag;
  wire       [15:0]   twiddle_factor_table_1_real;
  wire       [15:0]   twiddle_factor_table_1_imag;
  wire       [15:0]   twiddle_factor_table_2_real;
  wire       [15:0]   twiddle_factor_table_2_imag;
  wire       [15:0]   twiddle_factor_table_3_real;
  wire       [15:0]   twiddle_factor_table_3_imag;
  wire       [15:0]   twiddle_factor_table_4_real;
  wire       [15:0]   twiddle_factor_table_4_imag;
  wire       [15:0]   twiddle_factor_table_5_real;
  wire       [15:0]   twiddle_factor_table_5_imag;
  wire       [15:0]   twiddle_factor_table_6_real;
  wire       [15:0]   twiddle_factor_table_6_imag;
  wire       [15:0]   twiddle_factor_table_7_real;
  wire       [15:0]   twiddle_factor_table_7_imag;
  wire       [15:0]   twiddle_factor_table_8_real;
  wire       [15:0]   twiddle_factor_table_8_imag;
  wire       [15:0]   twiddle_factor_table_9_real;
  wire       [15:0]   twiddle_factor_table_9_imag;
  wire       [15:0]   twiddle_factor_table_10_real;
  wire       [15:0]   twiddle_factor_table_10_imag;
  wire       [15:0]   twiddle_factor_table_11_real;
  wire       [15:0]   twiddle_factor_table_11_imag;
  wire       [15:0]   twiddle_factor_table_12_real;
  wire       [15:0]   twiddle_factor_table_12_imag;
  wire       [15:0]   twiddle_factor_table_13_real;
  wire       [15:0]   twiddle_factor_table_13_imag;
  wire       [15:0]   twiddle_factor_table_14_real;
  wire       [15:0]   twiddle_factor_table_14_imag;
  wire       [15:0]   twiddle_factor_table_15_real;
  wire       [15:0]   twiddle_factor_table_15_imag;
  wire       [15:0]   twiddle_factor_table_16_real;
  wire       [15:0]   twiddle_factor_table_16_imag;
  wire       [15:0]   twiddle_factor_table_17_real;
  wire       [15:0]   twiddle_factor_table_17_imag;
  wire       [15:0]   twiddle_factor_table_18_real;
  wire       [15:0]   twiddle_factor_table_18_imag;
  wire       [15:0]   twiddle_factor_table_19_real;
  wire       [15:0]   twiddle_factor_table_19_imag;
  wire       [15:0]   twiddle_factor_table_20_real;
  wire       [15:0]   twiddle_factor_table_20_imag;
  wire       [15:0]   twiddle_factor_table_21_real;
  wire       [15:0]   twiddle_factor_table_21_imag;
  wire       [15:0]   twiddle_factor_table_22_real;
  wire       [15:0]   twiddle_factor_table_22_imag;
  wire       [15:0]   twiddle_factor_table_23_real;
  wire       [15:0]   twiddle_factor_table_23_imag;
  wire       [15:0]   twiddle_factor_table_24_real;
  wire       [15:0]   twiddle_factor_table_24_imag;
  wire       [15:0]   twiddle_factor_table_25_real;
  wire       [15:0]   twiddle_factor_table_25_imag;
  wire       [15:0]   twiddle_factor_table_26_real;
  wire       [15:0]   twiddle_factor_table_26_imag;
  wire       [15:0]   twiddle_factor_table_27_real;
  wire       [15:0]   twiddle_factor_table_27_imag;
  wire       [15:0]   twiddle_factor_table_28_real;
  wire       [15:0]   twiddle_factor_table_28_imag;
  wire       [15:0]   twiddle_factor_table_29_real;
  wire       [15:0]   twiddle_factor_table_29_imag;
  wire       [15:0]   twiddle_factor_table_30_real;
  wire       [15:0]   twiddle_factor_table_30_imag;
  wire       [15:0]   twiddle_factor_table_31_real;
  wire       [15:0]   twiddle_factor_table_31_imag;
  wire       [15:0]   twiddle_factor_table_32_real;
  wire       [15:0]   twiddle_factor_table_32_imag;
  wire       [15:0]   twiddle_factor_table_33_real;
  wire       [15:0]   twiddle_factor_table_33_imag;
  wire       [15:0]   twiddle_factor_table_34_real;
  wire       [15:0]   twiddle_factor_table_34_imag;
  wire       [15:0]   twiddle_factor_table_35_real;
  wire       [15:0]   twiddle_factor_table_35_imag;
  wire       [15:0]   twiddle_factor_table_36_real;
  wire       [15:0]   twiddle_factor_table_36_imag;
  wire       [15:0]   twiddle_factor_table_37_real;
  wire       [15:0]   twiddle_factor_table_37_imag;
  wire       [15:0]   twiddle_factor_table_38_real;
  wire       [15:0]   twiddle_factor_table_38_imag;
  wire       [15:0]   twiddle_factor_table_39_real;
  wire       [15:0]   twiddle_factor_table_39_imag;
  wire       [15:0]   twiddle_factor_table_40_real;
  wire       [15:0]   twiddle_factor_table_40_imag;
  wire       [15:0]   twiddle_factor_table_41_real;
  wire       [15:0]   twiddle_factor_table_41_imag;
  wire       [15:0]   twiddle_factor_table_42_real;
  wire       [15:0]   twiddle_factor_table_42_imag;
  wire       [15:0]   twiddle_factor_table_43_real;
  wire       [15:0]   twiddle_factor_table_43_imag;
  wire       [15:0]   twiddle_factor_table_44_real;
  wire       [15:0]   twiddle_factor_table_44_imag;
  wire       [15:0]   twiddle_factor_table_45_real;
  wire       [15:0]   twiddle_factor_table_45_imag;
  wire       [15:0]   twiddle_factor_table_46_real;
  wire       [15:0]   twiddle_factor_table_46_imag;
  wire       [15:0]   twiddle_factor_table_47_real;
  wire       [15:0]   twiddle_factor_table_47_imag;
  wire       [15:0]   twiddle_factor_table_48_real;
  wire       [15:0]   twiddle_factor_table_48_imag;
  wire       [15:0]   twiddle_factor_table_49_real;
  wire       [15:0]   twiddle_factor_table_49_imag;
  wire       [15:0]   twiddle_factor_table_50_real;
  wire       [15:0]   twiddle_factor_table_50_imag;
  wire       [15:0]   twiddle_factor_table_51_real;
  wire       [15:0]   twiddle_factor_table_51_imag;
  wire       [15:0]   twiddle_factor_table_52_real;
  wire       [15:0]   twiddle_factor_table_52_imag;
  wire       [15:0]   twiddle_factor_table_53_real;
  wire       [15:0]   twiddle_factor_table_53_imag;
  wire       [15:0]   twiddle_factor_table_54_real;
  wire       [15:0]   twiddle_factor_table_54_imag;
  wire       [15:0]   twiddle_factor_table_55_real;
  wire       [15:0]   twiddle_factor_table_55_imag;
  wire       [15:0]   twiddle_factor_table_56_real;
  wire       [15:0]   twiddle_factor_table_56_imag;
  wire       [15:0]   twiddle_factor_table_57_real;
  wire       [15:0]   twiddle_factor_table_57_imag;
  wire       [15:0]   twiddle_factor_table_58_real;
  wire       [15:0]   twiddle_factor_table_58_imag;
  wire       [15:0]   twiddle_factor_table_59_real;
  wire       [15:0]   twiddle_factor_table_59_imag;
  wire       [15:0]   twiddle_factor_table_60_real;
  wire       [15:0]   twiddle_factor_table_60_imag;
  wire       [15:0]   twiddle_factor_table_61_real;
  wire       [15:0]   twiddle_factor_table_61_imag;
  wire       [15:0]   twiddle_factor_table_62_real;
  wire       [15:0]   twiddle_factor_table_62_imag;
  wire       [15:0]   twiddle_factor_table_63_real;
  wire       [15:0]   twiddle_factor_table_63_imag;
  wire       [15:0]   twiddle_factor_table_64_real;
  wire       [15:0]   twiddle_factor_table_64_imag;
  wire       [15:0]   twiddle_factor_table_65_real;
  wire       [15:0]   twiddle_factor_table_65_imag;
  wire       [15:0]   twiddle_factor_table_66_real;
  wire       [15:0]   twiddle_factor_table_66_imag;
  wire       [15:0]   twiddle_factor_table_67_real;
  wire       [15:0]   twiddle_factor_table_67_imag;
  wire       [15:0]   twiddle_factor_table_68_real;
  wire       [15:0]   twiddle_factor_table_68_imag;
  wire       [15:0]   twiddle_factor_table_69_real;
  wire       [15:0]   twiddle_factor_table_69_imag;
  wire       [15:0]   twiddle_factor_table_70_real;
  wire       [15:0]   twiddle_factor_table_70_imag;
  wire       [15:0]   twiddle_factor_table_71_real;
  wire       [15:0]   twiddle_factor_table_71_imag;
  wire       [15:0]   twiddle_factor_table_72_real;
  wire       [15:0]   twiddle_factor_table_72_imag;
  wire       [15:0]   twiddle_factor_table_73_real;
  wire       [15:0]   twiddle_factor_table_73_imag;
  wire       [15:0]   twiddle_factor_table_74_real;
  wire       [15:0]   twiddle_factor_table_74_imag;
  wire       [15:0]   twiddle_factor_table_75_real;
  wire       [15:0]   twiddle_factor_table_75_imag;
  wire       [15:0]   twiddle_factor_table_76_real;
  wire       [15:0]   twiddle_factor_table_76_imag;
  wire       [15:0]   twiddle_factor_table_77_real;
  wire       [15:0]   twiddle_factor_table_77_imag;
  wire       [15:0]   twiddle_factor_table_78_real;
  wire       [15:0]   twiddle_factor_table_78_imag;
  wire       [15:0]   twiddle_factor_table_79_real;
  wire       [15:0]   twiddle_factor_table_79_imag;
  wire       [15:0]   twiddle_factor_table_80_real;
  wire       [15:0]   twiddle_factor_table_80_imag;
  wire       [15:0]   twiddle_factor_table_81_real;
  wire       [15:0]   twiddle_factor_table_81_imag;
  wire       [15:0]   twiddle_factor_table_82_real;
  wire       [15:0]   twiddle_factor_table_82_imag;
  wire       [15:0]   twiddle_factor_table_83_real;
  wire       [15:0]   twiddle_factor_table_83_imag;
  wire       [15:0]   twiddle_factor_table_84_real;
  wire       [15:0]   twiddle_factor_table_84_imag;
  wire       [15:0]   twiddle_factor_table_85_real;
  wire       [15:0]   twiddle_factor_table_85_imag;
  wire       [15:0]   twiddle_factor_table_86_real;
  wire       [15:0]   twiddle_factor_table_86_imag;
  wire       [15:0]   twiddle_factor_table_87_real;
  wire       [15:0]   twiddle_factor_table_87_imag;
  wire       [15:0]   twiddle_factor_table_88_real;
  wire       [15:0]   twiddle_factor_table_88_imag;
  wire       [15:0]   twiddle_factor_table_89_real;
  wire       [15:0]   twiddle_factor_table_89_imag;
  wire       [15:0]   twiddle_factor_table_90_real;
  wire       [15:0]   twiddle_factor_table_90_imag;
  wire       [15:0]   twiddle_factor_table_91_real;
  wire       [15:0]   twiddle_factor_table_91_imag;
  wire       [15:0]   twiddle_factor_table_92_real;
  wire       [15:0]   twiddle_factor_table_92_imag;
  wire       [15:0]   twiddle_factor_table_93_real;
  wire       [15:0]   twiddle_factor_table_93_imag;
  wire       [15:0]   twiddle_factor_table_94_real;
  wire       [15:0]   twiddle_factor_table_94_imag;
  wire       [15:0]   twiddle_factor_table_95_real;
  wire       [15:0]   twiddle_factor_table_95_imag;
  wire       [15:0]   twiddle_factor_table_96_real;
  wire       [15:0]   twiddle_factor_table_96_imag;
  wire       [15:0]   twiddle_factor_table_97_real;
  wire       [15:0]   twiddle_factor_table_97_imag;
  wire       [15:0]   twiddle_factor_table_98_real;
  wire       [15:0]   twiddle_factor_table_98_imag;
  wire       [15:0]   twiddle_factor_table_99_real;
  wire       [15:0]   twiddle_factor_table_99_imag;
  wire       [15:0]   twiddle_factor_table_100_real;
  wire       [15:0]   twiddle_factor_table_100_imag;
  wire       [15:0]   twiddle_factor_table_101_real;
  wire       [15:0]   twiddle_factor_table_101_imag;
  wire       [15:0]   twiddle_factor_table_102_real;
  wire       [15:0]   twiddle_factor_table_102_imag;
  wire       [15:0]   twiddle_factor_table_103_real;
  wire       [15:0]   twiddle_factor_table_103_imag;
  wire       [15:0]   twiddle_factor_table_104_real;
  wire       [15:0]   twiddle_factor_table_104_imag;
  wire       [15:0]   twiddle_factor_table_105_real;
  wire       [15:0]   twiddle_factor_table_105_imag;
  wire       [15:0]   twiddle_factor_table_106_real;
  wire       [15:0]   twiddle_factor_table_106_imag;
  wire       [15:0]   twiddle_factor_table_107_real;
  wire       [15:0]   twiddle_factor_table_107_imag;
  wire       [15:0]   twiddle_factor_table_108_real;
  wire       [15:0]   twiddle_factor_table_108_imag;
  wire       [15:0]   twiddle_factor_table_109_real;
  wire       [15:0]   twiddle_factor_table_109_imag;
  wire       [15:0]   twiddle_factor_table_110_real;
  wire       [15:0]   twiddle_factor_table_110_imag;
  wire       [15:0]   twiddle_factor_table_111_real;
  wire       [15:0]   twiddle_factor_table_111_imag;
  wire       [15:0]   twiddle_factor_table_112_real;
  wire       [15:0]   twiddle_factor_table_112_imag;
  wire       [15:0]   twiddle_factor_table_113_real;
  wire       [15:0]   twiddle_factor_table_113_imag;
  wire       [15:0]   twiddle_factor_table_114_real;
  wire       [15:0]   twiddle_factor_table_114_imag;
  wire       [15:0]   twiddle_factor_table_115_real;
  wire       [15:0]   twiddle_factor_table_115_imag;
  wire       [15:0]   twiddle_factor_table_116_real;
  wire       [15:0]   twiddle_factor_table_116_imag;
  wire       [15:0]   twiddle_factor_table_117_real;
  wire       [15:0]   twiddle_factor_table_117_imag;
  wire       [15:0]   twiddle_factor_table_118_real;
  wire       [15:0]   twiddle_factor_table_118_imag;
  wire       [15:0]   twiddle_factor_table_119_real;
  wire       [15:0]   twiddle_factor_table_119_imag;
  wire       [15:0]   twiddle_factor_table_120_real;
  wire       [15:0]   twiddle_factor_table_120_imag;
  wire       [15:0]   twiddle_factor_table_121_real;
  wire       [15:0]   twiddle_factor_table_121_imag;
  wire       [15:0]   twiddle_factor_table_122_real;
  wire       [15:0]   twiddle_factor_table_122_imag;
  wire       [15:0]   twiddle_factor_table_123_real;
  wire       [15:0]   twiddle_factor_table_123_imag;
  wire       [15:0]   twiddle_factor_table_124_real;
  wire       [15:0]   twiddle_factor_table_124_imag;
  wire       [15:0]   twiddle_factor_table_125_real;
  wire       [15:0]   twiddle_factor_table_125_imag;
  wire       [15:0]   twiddle_factor_table_126_real;
  wire       [15:0]   twiddle_factor_table_126_imag;
  wire       [15:0]   data_reorder_0_real;
  wire       [15:0]   data_reorder_0_imag;
  wire       [15:0]   data_reorder_1_real;
  wire       [15:0]   data_reorder_1_imag;
  wire       [15:0]   data_reorder_2_real;
  wire       [15:0]   data_reorder_2_imag;
  wire       [15:0]   data_reorder_3_real;
  wire       [15:0]   data_reorder_3_imag;
  wire       [15:0]   data_reorder_4_real;
  wire       [15:0]   data_reorder_4_imag;
  wire       [15:0]   data_reorder_5_real;
  wire       [15:0]   data_reorder_5_imag;
  wire       [15:0]   data_reorder_6_real;
  wire       [15:0]   data_reorder_6_imag;
  wire       [15:0]   data_reorder_7_real;
  wire       [15:0]   data_reorder_7_imag;
  wire       [15:0]   data_reorder_8_real;
  wire       [15:0]   data_reorder_8_imag;
  wire       [15:0]   data_reorder_9_real;
  wire       [15:0]   data_reorder_9_imag;
  wire       [15:0]   data_reorder_10_real;
  wire       [15:0]   data_reorder_10_imag;
  wire       [15:0]   data_reorder_11_real;
  wire       [15:0]   data_reorder_11_imag;
  wire       [15:0]   data_reorder_12_real;
  wire       [15:0]   data_reorder_12_imag;
  wire       [15:0]   data_reorder_13_real;
  wire       [15:0]   data_reorder_13_imag;
  wire       [15:0]   data_reorder_14_real;
  wire       [15:0]   data_reorder_14_imag;
  wire       [15:0]   data_reorder_15_real;
  wire       [15:0]   data_reorder_15_imag;
  wire       [15:0]   data_reorder_16_real;
  wire       [15:0]   data_reorder_16_imag;
  wire       [15:0]   data_reorder_17_real;
  wire       [15:0]   data_reorder_17_imag;
  wire       [15:0]   data_reorder_18_real;
  wire       [15:0]   data_reorder_18_imag;
  wire       [15:0]   data_reorder_19_real;
  wire       [15:0]   data_reorder_19_imag;
  wire       [15:0]   data_reorder_20_real;
  wire       [15:0]   data_reorder_20_imag;
  wire       [15:0]   data_reorder_21_real;
  wire       [15:0]   data_reorder_21_imag;
  wire       [15:0]   data_reorder_22_real;
  wire       [15:0]   data_reorder_22_imag;
  wire       [15:0]   data_reorder_23_real;
  wire       [15:0]   data_reorder_23_imag;
  wire       [15:0]   data_reorder_24_real;
  wire       [15:0]   data_reorder_24_imag;
  wire       [15:0]   data_reorder_25_real;
  wire       [15:0]   data_reorder_25_imag;
  wire       [15:0]   data_reorder_26_real;
  wire       [15:0]   data_reorder_26_imag;
  wire       [15:0]   data_reorder_27_real;
  wire       [15:0]   data_reorder_27_imag;
  wire       [15:0]   data_reorder_28_real;
  wire       [15:0]   data_reorder_28_imag;
  wire       [15:0]   data_reorder_29_real;
  wire       [15:0]   data_reorder_29_imag;
  wire       [15:0]   data_reorder_30_real;
  wire       [15:0]   data_reorder_30_imag;
  wire       [15:0]   data_reorder_31_real;
  wire       [15:0]   data_reorder_31_imag;
  wire       [15:0]   data_reorder_32_real;
  wire       [15:0]   data_reorder_32_imag;
  wire       [15:0]   data_reorder_33_real;
  wire       [15:0]   data_reorder_33_imag;
  wire       [15:0]   data_reorder_34_real;
  wire       [15:0]   data_reorder_34_imag;
  wire       [15:0]   data_reorder_35_real;
  wire       [15:0]   data_reorder_35_imag;
  wire       [15:0]   data_reorder_36_real;
  wire       [15:0]   data_reorder_36_imag;
  wire       [15:0]   data_reorder_37_real;
  wire       [15:0]   data_reorder_37_imag;
  wire       [15:0]   data_reorder_38_real;
  wire       [15:0]   data_reorder_38_imag;
  wire       [15:0]   data_reorder_39_real;
  wire       [15:0]   data_reorder_39_imag;
  wire       [15:0]   data_reorder_40_real;
  wire       [15:0]   data_reorder_40_imag;
  wire       [15:0]   data_reorder_41_real;
  wire       [15:0]   data_reorder_41_imag;
  wire       [15:0]   data_reorder_42_real;
  wire       [15:0]   data_reorder_42_imag;
  wire       [15:0]   data_reorder_43_real;
  wire       [15:0]   data_reorder_43_imag;
  wire       [15:0]   data_reorder_44_real;
  wire       [15:0]   data_reorder_44_imag;
  wire       [15:0]   data_reorder_45_real;
  wire       [15:0]   data_reorder_45_imag;
  wire       [15:0]   data_reorder_46_real;
  wire       [15:0]   data_reorder_46_imag;
  wire       [15:0]   data_reorder_47_real;
  wire       [15:0]   data_reorder_47_imag;
  wire       [15:0]   data_reorder_48_real;
  wire       [15:0]   data_reorder_48_imag;
  wire       [15:0]   data_reorder_49_real;
  wire       [15:0]   data_reorder_49_imag;
  wire       [15:0]   data_reorder_50_real;
  wire       [15:0]   data_reorder_50_imag;
  wire       [15:0]   data_reorder_51_real;
  wire       [15:0]   data_reorder_51_imag;
  wire       [15:0]   data_reorder_52_real;
  wire       [15:0]   data_reorder_52_imag;
  wire       [15:0]   data_reorder_53_real;
  wire       [15:0]   data_reorder_53_imag;
  wire       [15:0]   data_reorder_54_real;
  wire       [15:0]   data_reorder_54_imag;
  wire       [15:0]   data_reorder_55_real;
  wire       [15:0]   data_reorder_55_imag;
  wire       [15:0]   data_reorder_56_real;
  wire       [15:0]   data_reorder_56_imag;
  wire       [15:0]   data_reorder_57_real;
  wire       [15:0]   data_reorder_57_imag;
  wire       [15:0]   data_reorder_58_real;
  wire       [15:0]   data_reorder_58_imag;
  wire       [15:0]   data_reorder_59_real;
  wire       [15:0]   data_reorder_59_imag;
  wire       [15:0]   data_reorder_60_real;
  wire       [15:0]   data_reorder_60_imag;
  wire       [15:0]   data_reorder_61_real;
  wire       [15:0]   data_reorder_61_imag;
  wire       [15:0]   data_reorder_62_real;
  wire       [15:0]   data_reorder_62_imag;
  wire       [15:0]   data_reorder_63_real;
  wire       [15:0]   data_reorder_63_imag;
  wire       [15:0]   data_reorder_64_real;
  wire       [15:0]   data_reorder_64_imag;
  wire       [15:0]   data_reorder_65_real;
  wire       [15:0]   data_reorder_65_imag;
  wire       [15:0]   data_reorder_66_real;
  wire       [15:0]   data_reorder_66_imag;
  wire       [15:0]   data_reorder_67_real;
  wire       [15:0]   data_reorder_67_imag;
  wire       [15:0]   data_reorder_68_real;
  wire       [15:0]   data_reorder_68_imag;
  wire       [15:0]   data_reorder_69_real;
  wire       [15:0]   data_reorder_69_imag;
  wire       [15:0]   data_reorder_70_real;
  wire       [15:0]   data_reorder_70_imag;
  wire       [15:0]   data_reorder_71_real;
  wire       [15:0]   data_reorder_71_imag;
  wire       [15:0]   data_reorder_72_real;
  wire       [15:0]   data_reorder_72_imag;
  wire       [15:0]   data_reorder_73_real;
  wire       [15:0]   data_reorder_73_imag;
  wire       [15:0]   data_reorder_74_real;
  wire       [15:0]   data_reorder_74_imag;
  wire       [15:0]   data_reorder_75_real;
  wire       [15:0]   data_reorder_75_imag;
  wire       [15:0]   data_reorder_76_real;
  wire       [15:0]   data_reorder_76_imag;
  wire       [15:0]   data_reorder_77_real;
  wire       [15:0]   data_reorder_77_imag;
  wire       [15:0]   data_reorder_78_real;
  wire       [15:0]   data_reorder_78_imag;
  wire       [15:0]   data_reorder_79_real;
  wire       [15:0]   data_reorder_79_imag;
  wire       [15:0]   data_reorder_80_real;
  wire       [15:0]   data_reorder_80_imag;
  wire       [15:0]   data_reorder_81_real;
  wire       [15:0]   data_reorder_81_imag;
  wire       [15:0]   data_reorder_82_real;
  wire       [15:0]   data_reorder_82_imag;
  wire       [15:0]   data_reorder_83_real;
  wire       [15:0]   data_reorder_83_imag;
  wire       [15:0]   data_reorder_84_real;
  wire       [15:0]   data_reorder_84_imag;
  wire       [15:0]   data_reorder_85_real;
  wire       [15:0]   data_reorder_85_imag;
  wire       [15:0]   data_reorder_86_real;
  wire       [15:0]   data_reorder_86_imag;
  wire       [15:0]   data_reorder_87_real;
  wire       [15:0]   data_reorder_87_imag;
  wire       [15:0]   data_reorder_88_real;
  wire       [15:0]   data_reorder_88_imag;
  wire       [15:0]   data_reorder_89_real;
  wire       [15:0]   data_reorder_89_imag;
  wire       [15:0]   data_reorder_90_real;
  wire       [15:0]   data_reorder_90_imag;
  wire       [15:0]   data_reorder_91_real;
  wire       [15:0]   data_reorder_91_imag;
  wire       [15:0]   data_reorder_92_real;
  wire       [15:0]   data_reorder_92_imag;
  wire       [15:0]   data_reorder_93_real;
  wire       [15:0]   data_reorder_93_imag;
  wire       [15:0]   data_reorder_94_real;
  wire       [15:0]   data_reorder_94_imag;
  wire       [15:0]   data_reorder_95_real;
  wire       [15:0]   data_reorder_95_imag;
  wire       [15:0]   data_reorder_96_real;
  wire       [15:0]   data_reorder_96_imag;
  wire       [15:0]   data_reorder_97_real;
  wire       [15:0]   data_reorder_97_imag;
  wire       [15:0]   data_reorder_98_real;
  wire       [15:0]   data_reorder_98_imag;
  wire       [15:0]   data_reorder_99_real;
  wire       [15:0]   data_reorder_99_imag;
  wire       [15:0]   data_reorder_100_real;
  wire       [15:0]   data_reorder_100_imag;
  wire       [15:0]   data_reorder_101_real;
  wire       [15:0]   data_reorder_101_imag;
  wire       [15:0]   data_reorder_102_real;
  wire       [15:0]   data_reorder_102_imag;
  wire       [15:0]   data_reorder_103_real;
  wire       [15:0]   data_reorder_103_imag;
  wire       [15:0]   data_reorder_104_real;
  wire       [15:0]   data_reorder_104_imag;
  wire       [15:0]   data_reorder_105_real;
  wire       [15:0]   data_reorder_105_imag;
  wire       [15:0]   data_reorder_106_real;
  wire       [15:0]   data_reorder_106_imag;
  wire       [15:0]   data_reorder_107_real;
  wire       [15:0]   data_reorder_107_imag;
  wire       [15:0]   data_reorder_108_real;
  wire       [15:0]   data_reorder_108_imag;
  wire       [15:0]   data_reorder_109_real;
  wire       [15:0]   data_reorder_109_imag;
  wire       [15:0]   data_reorder_110_real;
  wire       [15:0]   data_reorder_110_imag;
  wire       [15:0]   data_reorder_111_real;
  wire       [15:0]   data_reorder_111_imag;
  wire       [15:0]   data_reorder_112_real;
  wire       [15:0]   data_reorder_112_imag;
  wire       [15:0]   data_reorder_113_real;
  wire       [15:0]   data_reorder_113_imag;
  wire       [15:0]   data_reorder_114_real;
  wire       [15:0]   data_reorder_114_imag;
  wire       [15:0]   data_reorder_115_real;
  wire       [15:0]   data_reorder_115_imag;
  wire       [15:0]   data_reorder_116_real;
  wire       [15:0]   data_reorder_116_imag;
  wire       [15:0]   data_reorder_117_real;
  wire       [15:0]   data_reorder_117_imag;
  wire       [15:0]   data_reorder_118_real;
  wire       [15:0]   data_reorder_118_imag;
  wire       [15:0]   data_reorder_119_real;
  wire       [15:0]   data_reorder_119_imag;
  wire       [15:0]   data_reorder_120_real;
  wire       [15:0]   data_reorder_120_imag;
  wire       [15:0]   data_reorder_121_real;
  wire       [15:0]   data_reorder_121_imag;
  wire       [15:0]   data_reorder_122_real;
  wire       [15:0]   data_reorder_122_imag;
  wire       [15:0]   data_reorder_123_real;
  wire       [15:0]   data_reorder_123_imag;
  wire       [15:0]   data_reorder_124_real;
  wire       [15:0]   data_reorder_124_imag;
  wire       [15:0]   data_reorder_125_real;
  wire       [15:0]   data_reorder_125_imag;
  wire       [15:0]   data_reorder_126_real;
  wire       [15:0]   data_reorder_126_imag;
  wire       [15:0]   data_reorder_127_real;
  wire       [15:0]   data_reorder_127_imag;
  reg        [15:0]   data_mid_0_real;
  reg        [15:0]   data_mid_0_imag;
  reg        [15:0]   data_mid_1_real;
  reg        [15:0]   data_mid_1_imag;
  reg        [15:0]   data_mid_2_real;
  reg        [15:0]   data_mid_2_imag;
  reg        [15:0]   data_mid_3_real;
  reg        [15:0]   data_mid_3_imag;
  reg        [15:0]   data_mid_4_real;
  reg        [15:0]   data_mid_4_imag;
  reg        [15:0]   data_mid_5_real;
  reg        [15:0]   data_mid_5_imag;
  reg        [15:0]   data_mid_6_real;
  reg        [15:0]   data_mid_6_imag;
  reg        [15:0]   data_mid_7_real;
  reg        [15:0]   data_mid_7_imag;
  reg        [15:0]   data_mid_8_real;
  reg        [15:0]   data_mid_8_imag;
  reg        [15:0]   data_mid_9_real;
  reg        [15:0]   data_mid_9_imag;
  reg        [15:0]   data_mid_10_real;
  reg        [15:0]   data_mid_10_imag;
  reg        [15:0]   data_mid_11_real;
  reg        [15:0]   data_mid_11_imag;
  reg        [15:0]   data_mid_12_real;
  reg        [15:0]   data_mid_12_imag;
  reg        [15:0]   data_mid_13_real;
  reg        [15:0]   data_mid_13_imag;
  reg        [15:0]   data_mid_14_real;
  reg        [15:0]   data_mid_14_imag;
  reg        [15:0]   data_mid_15_real;
  reg        [15:0]   data_mid_15_imag;
  reg        [15:0]   data_mid_16_real;
  reg        [15:0]   data_mid_16_imag;
  reg        [15:0]   data_mid_17_real;
  reg        [15:0]   data_mid_17_imag;
  reg        [15:0]   data_mid_18_real;
  reg        [15:0]   data_mid_18_imag;
  reg        [15:0]   data_mid_19_real;
  reg        [15:0]   data_mid_19_imag;
  reg        [15:0]   data_mid_20_real;
  reg        [15:0]   data_mid_20_imag;
  reg        [15:0]   data_mid_21_real;
  reg        [15:0]   data_mid_21_imag;
  reg        [15:0]   data_mid_22_real;
  reg        [15:0]   data_mid_22_imag;
  reg        [15:0]   data_mid_23_real;
  reg        [15:0]   data_mid_23_imag;
  reg        [15:0]   data_mid_24_real;
  reg        [15:0]   data_mid_24_imag;
  reg        [15:0]   data_mid_25_real;
  reg        [15:0]   data_mid_25_imag;
  reg        [15:0]   data_mid_26_real;
  reg        [15:0]   data_mid_26_imag;
  reg        [15:0]   data_mid_27_real;
  reg        [15:0]   data_mid_27_imag;
  reg        [15:0]   data_mid_28_real;
  reg        [15:0]   data_mid_28_imag;
  reg        [15:0]   data_mid_29_real;
  reg        [15:0]   data_mid_29_imag;
  reg        [15:0]   data_mid_30_real;
  reg        [15:0]   data_mid_30_imag;
  reg        [15:0]   data_mid_31_real;
  reg        [15:0]   data_mid_31_imag;
  reg        [15:0]   data_mid_32_real;
  reg        [15:0]   data_mid_32_imag;
  reg        [15:0]   data_mid_33_real;
  reg        [15:0]   data_mid_33_imag;
  reg        [15:0]   data_mid_34_real;
  reg        [15:0]   data_mid_34_imag;
  reg        [15:0]   data_mid_35_real;
  reg        [15:0]   data_mid_35_imag;
  reg        [15:0]   data_mid_36_real;
  reg        [15:0]   data_mid_36_imag;
  reg        [15:0]   data_mid_37_real;
  reg        [15:0]   data_mid_37_imag;
  reg        [15:0]   data_mid_38_real;
  reg        [15:0]   data_mid_38_imag;
  reg        [15:0]   data_mid_39_real;
  reg        [15:0]   data_mid_39_imag;
  reg        [15:0]   data_mid_40_real;
  reg        [15:0]   data_mid_40_imag;
  reg        [15:0]   data_mid_41_real;
  reg        [15:0]   data_mid_41_imag;
  reg        [15:0]   data_mid_42_real;
  reg        [15:0]   data_mid_42_imag;
  reg        [15:0]   data_mid_43_real;
  reg        [15:0]   data_mid_43_imag;
  reg        [15:0]   data_mid_44_real;
  reg        [15:0]   data_mid_44_imag;
  reg        [15:0]   data_mid_45_real;
  reg        [15:0]   data_mid_45_imag;
  reg        [15:0]   data_mid_46_real;
  reg        [15:0]   data_mid_46_imag;
  reg        [15:0]   data_mid_47_real;
  reg        [15:0]   data_mid_47_imag;
  reg        [15:0]   data_mid_48_real;
  reg        [15:0]   data_mid_48_imag;
  reg        [15:0]   data_mid_49_real;
  reg        [15:0]   data_mid_49_imag;
  reg        [15:0]   data_mid_50_real;
  reg        [15:0]   data_mid_50_imag;
  reg        [15:0]   data_mid_51_real;
  reg        [15:0]   data_mid_51_imag;
  reg        [15:0]   data_mid_52_real;
  reg        [15:0]   data_mid_52_imag;
  reg        [15:0]   data_mid_53_real;
  reg        [15:0]   data_mid_53_imag;
  reg        [15:0]   data_mid_54_real;
  reg        [15:0]   data_mid_54_imag;
  reg        [15:0]   data_mid_55_real;
  reg        [15:0]   data_mid_55_imag;
  reg        [15:0]   data_mid_56_real;
  reg        [15:0]   data_mid_56_imag;
  reg        [15:0]   data_mid_57_real;
  reg        [15:0]   data_mid_57_imag;
  reg        [15:0]   data_mid_58_real;
  reg        [15:0]   data_mid_58_imag;
  reg        [15:0]   data_mid_59_real;
  reg        [15:0]   data_mid_59_imag;
  reg        [15:0]   data_mid_60_real;
  reg        [15:0]   data_mid_60_imag;
  reg        [15:0]   data_mid_61_real;
  reg        [15:0]   data_mid_61_imag;
  reg        [15:0]   data_mid_62_real;
  reg        [15:0]   data_mid_62_imag;
  reg        [15:0]   data_mid_63_real;
  reg        [15:0]   data_mid_63_imag;
  reg        [15:0]   data_mid_64_real;
  reg        [15:0]   data_mid_64_imag;
  reg        [15:0]   data_mid_65_real;
  reg        [15:0]   data_mid_65_imag;
  reg        [15:0]   data_mid_66_real;
  reg        [15:0]   data_mid_66_imag;
  reg        [15:0]   data_mid_67_real;
  reg        [15:0]   data_mid_67_imag;
  reg        [15:0]   data_mid_68_real;
  reg        [15:0]   data_mid_68_imag;
  reg        [15:0]   data_mid_69_real;
  reg        [15:0]   data_mid_69_imag;
  reg        [15:0]   data_mid_70_real;
  reg        [15:0]   data_mid_70_imag;
  reg        [15:0]   data_mid_71_real;
  reg        [15:0]   data_mid_71_imag;
  reg        [15:0]   data_mid_72_real;
  reg        [15:0]   data_mid_72_imag;
  reg        [15:0]   data_mid_73_real;
  reg        [15:0]   data_mid_73_imag;
  reg        [15:0]   data_mid_74_real;
  reg        [15:0]   data_mid_74_imag;
  reg        [15:0]   data_mid_75_real;
  reg        [15:0]   data_mid_75_imag;
  reg        [15:0]   data_mid_76_real;
  reg        [15:0]   data_mid_76_imag;
  reg        [15:0]   data_mid_77_real;
  reg        [15:0]   data_mid_77_imag;
  reg        [15:0]   data_mid_78_real;
  reg        [15:0]   data_mid_78_imag;
  reg        [15:0]   data_mid_79_real;
  reg        [15:0]   data_mid_79_imag;
  reg        [15:0]   data_mid_80_real;
  reg        [15:0]   data_mid_80_imag;
  reg        [15:0]   data_mid_81_real;
  reg        [15:0]   data_mid_81_imag;
  reg        [15:0]   data_mid_82_real;
  reg        [15:0]   data_mid_82_imag;
  reg        [15:0]   data_mid_83_real;
  reg        [15:0]   data_mid_83_imag;
  reg        [15:0]   data_mid_84_real;
  reg        [15:0]   data_mid_84_imag;
  reg        [15:0]   data_mid_85_real;
  reg        [15:0]   data_mid_85_imag;
  reg        [15:0]   data_mid_86_real;
  reg        [15:0]   data_mid_86_imag;
  reg        [15:0]   data_mid_87_real;
  reg        [15:0]   data_mid_87_imag;
  reg        [15:0]   data_mid_88_real;
  reg        [15:0]   data_mid_88_imag;
  reg        [15:0]   data_mid_89_real;
  reg        [15:0]   data_mid_89_imag;
  reg        [15:0]   data_mid_90_real;
  reg        [15:0]   data_mid_90_imag;
  reg        [15:0]   data_mid_91_real;
  reg        [15:0]   data_mid_91_imag;
  reg        [15:0]   data_mid_92_real;
  reg        [15:0]   data_mid_92_imag;
  reg        [15:0]   data_mid_93_real;
  reg        [15:0]   data_mid_93_imag;
  reg        [15:0]   data_mid_94_real;
  reg        [15:0]   data_mid_94_imag;
  reg        [15:0]   data_mid_95_real;
  reg        [15:0]   data_mid_95_imag;
  reg        [15:0]   data_mid_96_real;
  reg        [15:0]   data_mid_96_imag;
  reg        [15:0]   data_mid_97_real;
  reg        [15:0]   data_mid_97_imag;
  reg        [15:0]   data_mid_98_real;
  reg        [15:0]   data_mid_98_imag;
  reg        [15:0]   data_mid_99_real;
  reg        [15:0]   data_mid_99_imag;
  reg        [15:0]   data_mid_100_real;
  reg        [15:0]   data_mid_100_imag;
  reg        [15:0]   data_mid_101_real;
  reg        [15:0]   data_mid_101_imag;
  reg        [15:0]   data_mid_102_real;
  reg        [15:0]   data_mid_102_imag;
  reg        [15:0]   data_mid_103_real;
  reg        [15:0]   data_mid_103_imag;
  reg        [15:0]   data_mid_104_real;
  reg        [15:0]   data_mid_104_imag;
  reg        [15:0]   data_mid_105_real;
  reg        [15:0]   data_mid_105_imag;
  reg        [15:0]   data_mid_106_real;
  reg        [15:0]   data_mid_106_imag;
  reg        [15:0]   data_mid_107_real;
  reg        [15:0]   data_mid_107_imag;
  reg        [15:0]   data_mid_108_real;
  reg        [15:0]   data_mid_108_imag;
  reg        [15:0]   data_mid_109_real;
  reg        [15:0]   data_mid_109_imag;
  reg        [15:0]   data_mid_110_real;
  reg        [15:0]   data_mid_110_imag;
  reg        [15:0]   data_mid_111_real;
  reg        [15:0]   data_mid_111_imag;
  reg        [15:0]   data_mid_112_real;
  reg        [15:0]   data_mid_112_imag;
  reg        [15:0]   data_mid_113_real;
  reg        [15:0]   data_mid_113_imag;
  reg        [15:0]   data_mid_114_real;
  reg        [15:0]   data_mid_114_imag;
  reg        [15:0]   data_mid_115_real;
  reg        [15:0]   data_mid_115_imag;
  reg        [15:0]   data_mid_116_real;
  reg        [15:0]   data_mid_116_imag;
  reg        [15:0]   data_mid_117_real;
  reg        [15:0]   data_mid_117_imag;
  reg        [15:0]   data_mid_118_real;
  reg        [15:0]   data_mid_118_imag;
  reg        [15:0]   data_mid_119_real;
  reg        [15:0]   data_mid_119_imag;
  reg        [15:0]   data_mid_120_real;
  reg        [15:0]   data_mid_120_imag;
  reg        [15:0]   data_mid_121_real;
  reg        [15:0]   data_mid_121_imag;
  reg        [15:0]   data_mid_122_real;
  reg        [15:0]   data_mid_122_imag;
  reg        [15:0]   data_mid_123_real;
  reg        [15:0]   data_mid_123_imag;
  reg        [15:0]   data_mid_124_real;
  reg        [15:0]   data_mid_124_imag;
  reg        [15:0]   data_mid_125_real;
  reg        [15:0]   data_mid_125_imag;
  reg        [15:0]   data_mid_126_real;
  reg        [15:0]   data_mid_126_imag;
  reg        [15:0]   data_mid_127_real;
  reg        [15:0]   data_mid_127_imag;
  reg                 io_data_in_valid_regNext;
  reg                 current_level_cnt_willIncrement;
  wire                current_level_cnt_willClear;
  reg        [2:0]    current_level_cnt_valueNext;
  reg        [2:0]    current_level_cnt_value;
  wire                current_level_cnt_willOverflowIfInc;
  wire                current_level_cnt_willOverflow;
  reg                 current_level_cond_period_minus_1;
  wire                current_level_cond_period;
  wire       [15:0]   _zz_1;
  wire       [15:0]   _zz_2;
  wire       [0:0]    _zz_3;
  wire       [0:0]    _zz_4;
  wire       [15:0]   _zz_5;
  wire       [15:0]   _zz_6;
  wire       [0:0]    _zz_7;
  wire       [0:0]    _zz_8;
  wire       [15:0]   _zz_9;
  wire       [15:0]   _zz_10;
  wire       [0:0]    _zz_11;
  wire       [0:0]    _zz_12;
  wire       [15:0]   _zz_13;
  wire       [15:0]   _zz_14;
  wire       [0:0]    _zz_15;
  wire       [0:0]    _zz_16;
  wire       [15:0]   _zz_17;
  wire       [15:0]   _zz_18;
  wire       [0:0]    _zz_19;
  wire       [0:0]    _zz_20;
  wire       [15:0]   _zz_21;
  wire       [15:0]   _zz_22;
  wire       [0:0]    _zz_23;
  wire       [0:0]    _zz_24;
  wire       [15:0]   _zz_25;
  wire       [15:0]   _zz_26;
  wire       [0:0]    _zz_27;
  wire       [0:0]    _zz_28;
  wire       [15:0]   _zz_29;
  wire       [15:0]   _zz_30;
  wire       [0:0]    _zz_31;
  wire       [0:0]    _zz_32;
  wire       [15:0]   _zz_33;
  wire       [15:0]   _zz_34;
  wire       [0:0]    _zz_35;
  wire       [0:0]    _zz_36;
  wire       [15:0]   _zz_37;
  wire       [15:0]   _zz_38;
  wire       [0:0]    _zz_39;
  wire       [0:0]    _zz_40;
  wire       [15:0]   _zz_41;
  wire       [15:0]   _zz_42;
  wire       [0:0]    _zz_43;
  wire       [0:0]    _zz_44;
  wire       [15:0]   _zz_45;
  wire       [15:0]   _zz_46;
  wire       [0:0]    _zz_47;
  wire       [0:0]    _zz_48;
  wire       [15:0]   _zz_49;
  wire       [15:0]   _zz_50;
  wire       [0:0]    _zz_51;
  wire       [0:0]    _zz_52;
  wire       [15:0]   _zz_53;
  wire       [15:0]   _zz_54;
  wire       [0:0]    _zz_55;
  wire       [0:0]    _zz_56;
  wire       [15:0]   _zz_57;
  wire       [15:0]   _zz_58;
  wire       [0:0]    _zz_59;
  wire       [0:0]    _zz_60;
  wire       [15:0]   _zz_61;
  wire       [15:0]   _zz_62;
  wire       [0:0]    _zz_63;
  wire       [0:0]    _zz_64;
  wire       [15:0]   _zz_65;
  wire       [15:0]   _zz_66;
  wire       [0:0]    _zz_67;
  wire       [0:0]    _zz_68;
  wire       [15:0]   _zz_69;
  wire       [15:0]   _zz_70;
  wire       [0:0]    _zz_71;
  wire       [0:0]    _zz_72;
  wire       [15:0]   _zz_73;
  wire       [15:0]   _zz_74;
  wire       [0:0]    _zz_75;
  wire       [0:0]    _zz_76;
  wire       [15:0]   _zz_77;
  wire       [15:0]   _zz_78;
  wire       [0:0]    _zz_79;
  wire       [0:0]    _zz_80;
  wire       [15:0]   _zz_81;
  wire       [15:0]   _zz_82;
  wire       [0:0]    _zz_83;
  wire       [0:0]    _zz_84;
  wire       [15:0]   _zz_85;
  wire       [15:0]   _zz_86;
  wire       [0:0]    _zz_87;
  wire       [0:0]    _zz_88;
  wire       [15:0]   _zz_89;
  wire       [15:0]   _zz_90;
  wire       [0:0]    _zz_91;
  wire       [0:0]    _zz_92;
  wire       [15:0]   _zz_93;
  wire       [15:0]   _zz_94;
  wire       [0:0]    _zz_95;
  wire       [0:0]    _zz_96;
  wire       [15:0]   _zz_97;
  wire       [15:0]   _zz_98;
  wire       [0:0]    _zz_99;
  wire       [0:0]    _zz_100;
  wire       [15:0]   _zz_101;
  wire       [15:0]   _zz_102;
  wire       [0:0]    _zz_103;
  wire       [0:0]    _zz_104;
  wire       [15:0]   _zz_105;
  wire       [15:0]   _zz_106;
  wire       [0:0]    _zz_107;
  wire       [0:0]    _zz_108;
  wire       [15:0]   _zz_109;
  wire       [15:0]   _zz_110;
  wire       [0:0]    _zz_111;
  wire       [0:0]    _zz_112;
  wire       [15:0]   _zz_113;
  wire       [15:0]   _zz_114;
  wire       [0:0]    _zz_115;
  wire       [0:0]    _zz_116;
  wire       [15:0]   _zz_117;
  wire       [15:0]   _zz_118;
  wire       [0:0]    _zz_119;
  wire       [0:0]    _zz_120;
  wire       [15:0]   _zz_121;
  wire       [15:0]   _zz_122;
  wire       [0:0]    _zz_123;
  wire       [0:0]    _zz_124;
  wire       [15:0]   _zz_125;
  wire       [15:0]   _zz_126;
  wire       [0:0]    _zz_127;
  wire       [0:0]    _zz_128;
  wire       [15:0]   _zz_129;
  wire       [15:0]   _zz_130;
  wire       [0:0]    _zz_131;
  wire       [0:0]    _zz_132;
  wire       [15:0]   _zz_133;
  wire       [15:0]   _zz_134;
  wire       [0:0]    _zz_135;
  wire       [0:0]    _zz_136;
  wire       [15:0]   _zz_137;
  wire       [15:0]   _zz_138;
  wire       [0:0]    _zz_139;
  wire       [0:0]    _zz_140;
  wire       [15:0]   _zz_141;
  wire       [15:0]   _zz_142;
  wire       [0:0]    _zz_143;
  wire       [0:0]    _zz_144;
  wire       [15:0]   _zz_145;
  wire       [15:0]   _zz_146;
  wire       [0:0]    _zz_147;
  wire       [0:0]    _zz_148;
  wire       [15:0]   _zz_149;
  wire       [15:0]   _zz_150;
  wire       [0:0]    _zz_151;
  wire       [0:0]    _zz_152;
  wire       [15:0]   _zz_153;
  wire       [15:0]   _zz_154;
  wire       [0:0]    _zz_155;
  wire       [0:0]    _zz_156;
  wire       [15:0]   _zz_157;
  wire       [15:0]   _zz_158;
  wire       [0:0]    _zz_159;
  wire       [0:0]    _zz_160;
  wire       [15:0]   _zz_161;
  wire       [15:0]   _zz_162;
  wire       [0:0]    _zz_163;
  wire       [0:0]    _zz_164;
  wire       [15:0]   _zz_165;
  wire       [15:0]   _zz_166;
  wire       [0:0]    _zz_167;
  wire       [0:0]    _zz_168;
  wire       [15:0]   _zz_169;
  wire       [15:0]   _zz_170;
  wire       [0:0]    _zz_171;
  wire       [0:0]    _zz_172;
  wire       [15:0]   _zz_173;
  wire       [15:0]   _zz_174;
  wire       [0:0]    _zz_175;
  wire       [0:0]    _zz_176;
  wire       [15:0]   _zz_177;
  wire       [15:0]   _zz_178;
  wire       [0:0]    _zz_179;
  wire       [0:0]    _zz_180;
  wire       [15:0]   _zz_181;
  wire       [15:0]   _zz_182;
  wire       [0:0]    _zz_183;
  wire       [0:0]    _zz_184;
  wire       [15:0]   _zz_185;
  wire       [15:0]   _zz_186;
  wire       [0:0]    _zz_187;
  wire       [0:0]    _zz_188;
  wire       [15:0]   _zz_189;
  wire       [15:0]   _zz_190;
  wire       [0:0]    _zz_191;
  wire       [0:0]    _zz_192;
  wire       [15:0]   _zz_193;
  wire       [15:0]   _zz_194;
  wire       [0:0]    _zz_195;
  wire       [0:0]    _zz_196;
  wire       [15:0]   _zz_197;
  wire       [15:0]   _zz_198;
  wire       [0:0]    _zz_199;
  wire       [0:0]    _zz_200;
  wire       [15:0]   _zz_201;
  wire       [15:0]   _zz_202;
  wire       [0:0]    _zz_203;
  wire       [0:0]    _zz_204;
  wire       [15:0]   _zz_205;
  wire       [15:0]   _zz_206;
  wire       [0:0]    _zz_207;
  wire       [0:0]    _zz_208;
  wire       [15:0]   _zz_209;
  wire       [15:0]   _zz_210;
  wire       [0:0]    _zz_211;
  wire       [0:0]    _zz_212;
  wire       [15:0]   _zz_213;
  wire       [15:0]   _zz_214;
  wire       [0:0]    _zz_215;
  wire       [0:0]    _zz_216;
  wire       [15:0]   _zz_217;
  wire       [15:0]   _zz_218;
  wire       [0:0]    _zz_219;
  wire       [0:0]    _zz_220;
  wire       [15:0]   _zz_221;
  wire       [15:0]   _zz_222;
  wire       [0:0]    _zz_223;
  wire       [0:0]    _zz_224;
  wire       [15:0]   _zz_225;
  wire       [15:0]   _zz_226;
  wire       [0:0]    _zz_227;
  wire       [0:0]    _zz_228;
  wire       [15:0]   _zz_229;
  wire       [15:0]   _zz_230;
  wire       [0:0]    _zz_231;
  wire       [0:0]    _zz_232;
  wire       [15:0]   _zz_233;
  wire       [15:0]   _zz_234;
  wire       [0:0]    _zz_235;
  wire       [0:0]    _zz_236;
  wire       [15:0]   _zz_237;
  wire       [15:0]   _zz_238;
  wire       [0:0]    _zz_239;
  wire       [0:0]    _zz_240;
  wire       [15:0]   _zz_241;
  wire       [15:0]   _zz_242;
  wire       [0:0]    _zz_243;
  wire       [0:0]    _zz_244;
  wire       [15:0]   _zz_245;
  wire       [15:0]   _zz_246;
  wire       [0:0]    _zz_247;
  wire       [0:0]    _zz_248;
  wire       [15:0]   _zz_249;
  wire       [15:0]   _zz_250;
  wire       [0:0]    _zz_251;
  wire       [0:0]    _zz_252;
  wire       [15:0]   _zz_253;
  wire       [15:0]   _zz_254;
  wire       [0:0]    _zz_255;
  wire       [0:0]    _zz_256;
  wire       [15:0]   _zz_257;
  wire       [15:0]   _zz_258;
  wire       [0:0]    _zz_259;
  wire       [0:0]    _zz_260;
  wire       [15:0]   _zz_261;
  wire       [15:0]   _zz_262;
  wire       [0:0]    _zz_263;
  wire       [0:0]    _zz_264;
  wire       [15:0]   _zz_265;
  wire       [15:0]   _zz_266;
  wire       [0:0]    _zz_267;
  wire       [0:0]    _zz_268;
  wire       [15:0]   _zz_269;
  wire       [15:0]   _zz_270;
  wire       [0:0]    _zz_271;
  wire       [0:0]    _zz_272;
  wire       [15:0]   _zz_273;
  wire       [15:0]   _zz_274;
  wire       [0:0]    _zz_275;
  wire       [0:0]    _zz_276;
  wire       [15:0]   _zz_277;
  wire       [15:0]   _zz_278;
  wire       [0:0]    _zz_279;
  wire       [0:0]    _zz_280;
  wire       [15:0]   _zz_281;
  wire       [15:0]   _zz_282;
  wire       [0:0]    _zz_283;
  wire       [0:0]    _zz_284;
  wire       [15:0]   _zz_285;
  wire       [15:0]   _zz_286;
  wire       [0:0]    _zz_287;
  wire       [0:0]    _zz_288;
  wire       [15:0]   _zz_289;
  wire       [15:0]   _zz_290;
  wire       [0:0]    _zz_291;
  wire       [0:0]    _zz_292;
  wire       [15:0]   _zz_293;
  wire       [15:0]   _zz_294;
  wire       [0:0]    _zz_295;
  wire       [0:0]    _zz_296;
  wire       [15:0]   _zz_297;
  wire       [15:0]   _zz_298;
  wire       [0:0]    _zz_299;
  wire       [0:0]    _zz_300;
  wire       [15:0]   _zz_301;
  wire       [15:0]   _zz_302;
  wire       [0:0]    _zz_303;
  wire       [0:0]    _zz_304;
  wire       [15:0]   _zz_305;
  wire       [15:0]   _zz_306;
  wire       [0:0]    _zz_307;
  wire       [0:0]    _zz_308;
  wire       [15:0]   _zz_309;
  wire       [15:0]   _zz_310;
  wire       [0:0]    _zz_311;
  wire       [0:0]    _zz_312;
  wire       [15:0]   _zz_313;
  wire       [15:0]   _zz_314;
  wire       [0:0]    _zz_315;
  wire       [0:0]    _zz_316;
  wire       [15:0]   _zz_317;
  wire       [15:0]   _zz_318;
  wire       [0:0]    _zz_319;
  wire       [0:0]    _zz_320;
  wire       [15:0]   _zz_321;
  wire       [15:0]   _zz_322;
  wire       [0:0]    _zz_323;
  wire       [0:0]    _zz_324;
  wire       [15:0]   _zz_325;
  wire       [15:0]   _zz_326;
  wire       [0:0]    _zz_327;
  wire       [0:0]    _zz_328;
  wire       [15:0]   _zz_329;
  wire       [15:0]   _zz_330;
  wire       [0:0]    _zz_331;
  wire       [0:0]    _zz_332;
  wire       [15:0]   _zz_333;
  wire       [15:0]   _zz_334;
  wire       [0:0]    _zz_335;
  wire       [0:0]    _zz_336;
  wire       [15:0]   _zz_337;
  wire       [15:0]   _zz_338;
  wire       [0:0]    _zz_339;
  wire       [0:0]    _zz_340;
  wire       [15:0]   _zz_341;
  wire       [15:0]   _zz_342;
  wire       [0:0]    _zz_343;
  wire       [0:0]    _zz_344;
  wire       [15:0]   _zz_345;
  wire       [15:0]   _zz_346;
  wire       [0:0]    _zz_347;
  wire       [0:0]    _zz_348;
  wire       [15:0]   _zz_349;
  wire       [15:0]   _zz_350;
  wire       [0:0]    _zz_351;
  wire       [0:0]    _zz_352;
  wire       [15:0]   _zz_353;
  wire       [15:0]   _zz_354;
  wire       [0:0]    _zz_355;
  wire       [0:0]    _zz_356;
  wire       [15:0]   _zz_357;
  wire       [15:0]   _zz_358;
  wire       [0:0]    _zz_359;
  wire       [0:0]    _zz_360;
  wire       [15:0]   _zz_361;
  wire       [15:0]   _zz_362;
  wire       [0:0]    _zz_363;
  wire       [0:0]    _zz_364;
  wire       [15:0]   _zz_365;
  wire       [15:0]   _zz_366;
  wire       [0:0]    _zz_367;
  wire       [0:0]    _zz_368;
  wire       [15:0]   _zz_369;
  wire       [15:0]   _zz_370;
  wire       [0:0]    _zz_371;
  wire       [0:0]    _zz_372;
  wire       [15:0]   _zz_373;
  wire       [15:0]   _zz_374;
  wire       [0:0]    _zz_375;
  wire       [0:0]    _zz_376;
  wire       [15:0]   _zz_377;
  wire       [15:0]   _zz_378;
  wire       [0:0]    _zz_379;
  wire       [0:0]    _zz_380;
  wire       [15:0]   _zz_381;
  wire       [15:0]   _zz_382;
  wire       [0:0]    _zz_383;
  wire       [0:0]    _zz_384;
  wire       [15:0]   _zz_385;
  wire       [15:0]   _zz_386;
  wire       [0:0]    _zz_387;
  wire       [0:0]    _zz_388;
  wire       [15:0]   _zz_389;
  wire       [15:0]   _zz_390;
  wire       [0:0]    _zz_391;
  wire       [0:0]    _zz_392;
  wire       [15:0]   _zz_393;
  wire       [15:0]   _zz_394;
  wire       [0:0]    _zz_395;
  wire       [0:0]    _zz_396;
  wire       [15:0]   _zz_397;
  wire       [15:0]   _zz_398;
  wire       [0:0]    _zz_399;
  wire       [0:0]    _zz_400;
  wire       [15:0]   _zz_401;
  wire       [15:0]   _zz_402;
  wire       [0:0]    _zz_403;
  wire       [0:0]    _zz_404;
  wire       [15:0]   _zz_405;
  wire       [15:0]   _zz_406;
  wire       [0:0]    _zz_407;
  wire       [0:0]    _zz_408;
  wire       [15:0]   _zz_409;
  wire       [15:0]   _zz_410;
  wire       [0:0]    _zz_411;
  wire       [0:0]    _zz_412;
  wire       [15:0]   _zz_413;
  wire       [15:0]   _zz_414;
  wire       [0:0]    _zz_415;
  wire       [0:0]    _zz_416;
  wire       [15:0]   _zz_417;
  wire       [15:0]   _zz_418;
  wire       [0:0]    _zz_419;
  wire       [0:0]    _zz_420;
  wire       [15:0]   _zz_421;
  wire       [15:0]   _zz_422;
  wire       [0:0]    _zz_423;
  wire       [0:0]    _zz_424;
  wire       [15:0]   _zz_425;
  wire       [15:0]   _zz_426;
  wire       [0:0]    _zz_427;
  wire       [0:0]    _zz_428;
  wire       [15:0]   _zz_429;
  wire       [15:0]   _zz_430;
  wire       [0:0]    _zz_431;
  wire       [0:0]    _zz_432;
  wire       [15:0]   _zz_433;
  wire       [15:0]   _zz_434;
  wire       [0:0]    _zz_435;
  wire       [0:0]    _zz_436;
  wire       [15:0]   _zz_437;
  wire       [15:0]   _zz_438;
  wire       [0:0]    _zz_439;
  wire       [0:0]    _zz_440;
  wire       [15:0]   _zz_441;
  wire       [15:0]   _zz_442;
  wire       [0:0]    _zz_443;
  wire       [0:0]    _zz_444;
  wire       [15:0]   _zz_445;
  wire       [15:0]   _zz_446;
  wire       [0:0]    _zz_447;
  wire       [0:0]    _zz_448;
  wire       [15:0]   _zz_449;
  wire       [15:0]   _zz_450;
  wire       [0:0]    _zz_451;
  wire       [0:0]    _zz_452;
  wire       [15:0]   _zz_453;
  wire       [15:0]   _zz_454;
  wire       [0:0]    _zz_455;
  wire       [0:0]    _zz_456;
  wire       [15:0]   _zz_457;
  wire       [15:0]   _zz_458;
  wire       [0:0]    _zz_459;
  wire       [0:0]    _zz_460;
  wire       [15:0]   _zz_461;
  wire       [15:0]   _zz_462;
  wire       [0:0]    _zz_463;
  wire       [0:0]    _zz_464;
  wire       [15:0]   _zz_465;
  wire       [15:0]   _zz_466;
  wire       [0:0]    _zz_467;
  wire       [0:0]    _zz_468;
  wire       [15:0]   _zz_469;
  wire       [15:0]   _zz_470;
  wire       [0:0]    _zz_471;
  wire       [0:0]    _zz_472;
  wire       [15:0]   _zz_473;
  wire       [15:0]   _zz_474;
  wire       [0:0]    _zz_475;
  wire       [0:0]    _zz_476;
  wire       [15:0]   _zz_477;
  wire       [15:0]   _zz_478;
  wire       [0:0]    _zz_479;
  wire       [0:0]    _zz_480;
  wire       [15:0]   _zz_481;
  wire       [15:0]   _zz_482;
  wire       [0:0]    _zz_483;
  wire       [0:0]    _zz_484;
  wire       [15:0]   _zz_485;
  wire       [15:0]   _zz_486;
  wire       [0:0]    _zz_487;
  wire       [0:0]    _zz_488;
  wire       [15:0]   _zz_489;
  wire       [15:0]   _zz_490;
  wire       [0:0]    _zz_491;
  wire       [0:0]    _zz_492;
  wire       [15:0]   _zz_493;
  wire       [15:0]   _zz_494;
  wire       [0:0]    _zz_495;
  wire       [0:0]    _zz_496;
  wire       [15:0]   _zz_497;
  wire       [15:0]   _zz_498;
  wire       [0:0]    _zz_499;
  wire       [0:0]    _zz_500;
  wire       [15:0]   _zz_501;
  wire       [15:0]   _zz_502;
  wire       [0:0]    _zz_503;
  wire       [0:0]    _zz_504;
  wire       [15:0]   _zz_505;
  wire       [15:0]   _zz_506;
  wire       [0:0]    _zz_507;
  wire       [0:0]    _zz_508;
  wire       [15:0]   _zz_509;
  wire       [15:0]   _zz_510;
  wire       [0:0]    _zz_511;
  wire       [0:0]    _zz_512;
  wire       [15:0]   _zz_513;
  wire       [15:0]   _zz_514;
  wire       [0:0]    _zz_515;
  wire       [0:0]    _zz_516;
  wire       [15:0]   _zz_517;
  wire       [15:0]   _zz_518;
  wire       [0:0]    _zz_519;
  wire       [0:0]    _zz_520;
  wire       [15:0]   _zz_521;
  wire       [15:0]   _zz_522;
  wire       [0:0]    _zz_523;
  wire       [0:0]    _zz_524;
  wire       [15:0]   _zz_525;
  wire       [15:0]   _zz_526;
  wire       [0:0]    _zz_527;
  wire       [0:0]    _zz_528;
  wire       [15:0]   _zz_529;
  wire       [15:0]   _zz_530;
  wire       [0:0]    _zz_531;
  wire       [0:0]    _zz_532;
  wire       [15:0]   _zz_533;
  wire       [15:0]   _zz_534;
  wire       [0:0]    _zz_535;
  wire       [0:0]    _zz_536;
  wire       [15:0]   _zz_537;
  wire       [15:0]   _zz_538;
  wire       [0:0]    _zz_539;
  wire       [0:0]    _zz_540;
  wire       [15:0]   _zz_541;
  wire       [15:0]   _zz_542;
  wire       [0:0]    _zz_543;
  wire       [0:0]    _zz_544;
  wire       [15:0]   _zz_545;
  wire       [15:0]   _zz_546;
  wire       [0:0]    _zz_547;
  wire       [0:0]    _zz_548;
  wire       [15:0]   _zz_549;
  wire       [15:0]   _zz_550;
  wire       [0:0]    _zz_551;
  wire       [0:0]    _zz_552;
  wire       [15:0]   _zz_553;
  wire       [15:0]   _zz_554;
  wire       [0:0]    _zz_555;
  wire       [0:0]    _zz_556;
  wire       [15:0]   _zz_557;
  wire       [15:0]   _zz_558;
  wire       [0:0]    _zz_559;
  wire       [0:0]    _zz_560;
  wire       [15:0]   _zz_561;
  wire       [15:0]   _zz_562;
  wire       [0:0]    _zz_563;
  wire       [0:0]    _zz_564;
  wire       [15:0]   _zz_565;
  wire       [15:0]   _zz_566;
  wire       [0:0]    _zz_567;
  wire       [0:0]    _zz_568;
  wire       [15:0]   _zz_569;
  wire       [15:0]   _zz_570;
  wire       [0:0]    _zz_571;
  wire       [0:0]    _zz_572;
  wire       [15:0]   _zz_573;
  wire       [15:0]   _zz_574;
  wire       [0:0]    _zz_575;
  wire       [0:0]    _zz_576;
  wire       [15:0]   _zz_577;
  wire       [15:0]   _zz_578;
  wire       [0:0]    _zz_579;
  wire       [0:0]    _zz_580;
  wire       [15:0]   _zz_581;
  wire       [15:0]   _zz_582;
  wire       [0:0]    _zz_583;
  wire       [0:0]    _zz_584;
  wire       [15:0]   _zz_585;
  wire       [15:0]   _zz_586;
  wire       [0:0]    _zz_587;
  wire       [0:0]    _zz_588;
  wire       [15:0]   _zz_589;
  wire       [15:0]   _zz_590;
  wire       [0:0]    _zz_591;
  wire       [0:0]    _zz_592;
  wire       [15:0]   _zz_593;
  wire       [15:0]   _zz_594;
  wire       [0:0]    _zz_595;
  wire       [0:0]    _zz_596;
  wire       [15:0]   _zz_597;
  wire       [15:0]   _zz_598;
  wire       [0:0]    _zz_599;
  wire       [0:0]    _zz_600;
  wire       [15:0]   _zz_601;
  wire       [15:0]   _zz_602;
  wire       [0:0]    _zz_603;
  wire       [0:0]    _zz_604;
  wire       [15:0]   _zz_605;
  wire       [15:0]   _zz_606;
  wire       [0:0]    _zz_607;
  wire       [0:0]    _zz_608;
  wire       [15:0]   _zz_609;
  wire       [15:0]   _zz_610;
  wire       [0:0]    _zz_611;
  wire       [0:0]    _zz_612;
  wire       [15:0]   _zz_613;
  wire       [15:0]   _zz_614;
  wire       [0:0]    _zz_615;
  wire       [0:0]    _zz_616;
  wire       [15:0]   _zz_617;
  wire       [15:0]   _zz_618;
  wire       [0:0]    _zz_619;
  wire       [0:0]    _zz_620;
  wire       [15:0]   _zz_621;
  wire       [15:0]   _zz_622;
  wire       [0:0]    _zz_623;
  wire       [0:0]    _zz_624;
  wire       [15:0]   _zz_625;
  wire       [15:0]   _zz_626;
  wire       [0:0]    _zz_627;
  wire       [0:0]    _zz_628;
  wire       [15:0]   _zz_629;
  wire       [15:0]   _zz_630;
  wire       [0:0]    _zz_631;
  wire       [0:0]    _zz_632;
  wire       [15:0]   _zz_633;
  wire       [15:0]   _zz_634;
  wire       [0:0]    _zz_635;
  wire       [0:0]    _zz_636;
  wire       [15:0]   _zz_637;
  wire       [15:0]   _zz_638;
  wire       [0:0]    _zz_639;
  wire       [0:0]    _zz_640;
  wire       [15:0]   _zz_641;
  wire       [15:0]   _zz_642;
  wire       [0:0]    _zz_643;
  wire       [0:0]    _zz_644;
  wire       [15:0]   _zz_645;
  wire       [15:0]   _zz_646;
  wire       [0:0]    _zz_647;
  wire       [0:0]    _zz_648;
  wire       [15:0]   _zz_649;
  wire       [15:0]   _zz_650;
  wire       [0:0]    _zz_651;
  wire       [0:0]    _zz_652;
  wire       [15:0]   _zz_653;
  wire       [15:0]   _zz_654;
  wire       [0:0]    _zz_655;
  wire       [0:0]    _zz_656;
  wire       [15:0]   _zz_657;
  wire       [15:0]   _zz_658;
  wire       [0:0]    _zz_659;
  wire       [0:0]    _zz_660;
  wire       [15:0]   _zz_661;
  wire       [15:0]   _zz_662;
  wire       [0:0]    _zz_663;
  wire       [0:0]    _zz_664;
  wire       [15:0]   _zz_665;
  wire       [15:0]   _zz_666;
  wire       [0:0]    _zz_667;
  wire       [0:0]    _zz_668;
  wire       [15:0]   _zz_669;
  wire       [15:0]   _zz_670;
  wire       [0:0]    _zz_671;
  wire       [0:0]    _zz_672;
  wire       [15:0]   _zz_673;
  wire       [15:0]   _zz_674;
  wire       [0:0]    _zz_675;
  wire       [0:0]    _zz_676;
  wire       [15:0]   _zz_677;
  wire       [15:0]   _zz_678;
  wire       [0:0]    _zz_679;
  wire       [0:0]    _zz_680;
  wire       [15:0]   _zz_681;
  wire       [15:0]   _zz_682;
  wire       [0:0]    _zz_683;
  wire       [0:0]    _zz_684;
  wire       [15:0]   _zz_685;
  wire       [15:0]   _zz_686;
  wire       [0:0]    _zz_687;
  wire       [0:0]    _zz_688;
  wire       [15:0]   _zz_689;
  wire       [15:0]   _zz_690;
  wire       [0:0]    _zz_691;
  wire       [0:0]    _zz_692;
  wire       [15:0]   _zz_693;
  wire       [15:0]   _zz_694;
  wire       [0:0]    _zz_695;
  wire       [0:0]    _zz_696;
  wire       [15:0]   _zz_697;
  wire       [15:0]   _zz_698;
  wire       [0:0]    _zz_699;
  wire       [0:0]    _zz_700;
  wire       [15:0]   _zz_701;
  wire       [15:0]   _zz_702;
  wire       [0:0]    _zz_703;
  wire       [0:0]    _zz_704;
  wire       [15:0]   _zz_705;
  wire       [15:0]   _zz_706;
  wire       [0:0]    _zz_707;
  wire       [0:0]    _zz_708;
  wire       [15:0]   _zz_709;
  wire       [15:0]   _zz_710;
  wire       [0:0]    _zz_711;
  wire       [0:0]    _zz_712;
  wire       [15:0]   _zz_713;
  wire       [15:0]   _zz_714;
  wire       [0:0]    _zz_715;
  wire       [0:0]    _zz_716;
  wire       [15:0]   _zz_717;
  wire       [15:0]   _zz_718;
  wire       [0:0]    _zz_719;
  wire       [0:0]    _zz_720;
  wire       [15:0]   _zz_721;
  wire       [15:0]   _zz_722;
  wire       [0:0]    _zz_723;
  wire       [0:0]    _zz_724;
  wire       [15:0]   _zz_725;
  wire       [15:0]   _zz_726;
  wire       [0:0]    _zz_727;
  wire       [0:0]    _zz_728;
  wire       [15:0]   _zz_729;
  wire       [15:0]   _zz_730;
  wire       [0:0]    _zz_731;
  wire       [0:0]    _zz_732;
  wire       [15:0]   _zz_733;
  wire       [15:0]   _zz_734;
  wire       [0:0]    _zz_735;
  wire       [0:0]    _zz_736;
  wire       [15:0]   _zz_737;
  wire       [15:0]   _zz_738;
  wire       [0:0]    _zz_739;
  wire       [0:0]    _zz_740;
  wire       [15:0]   _zz_741;
  wire       [15:0]   _zz_742;
  wire       [0:0]    _zz_743;
  wire       [0:0]    _zz_744;
  wire       [15:0]   _zz_745;
  wire       [15:0]   _zz_746;
  wire       [0:0]    _zz_747;
  wire       [0:0]    _zz_748;
  wire       [15:0]   _zz_749;
  wire       [15:0]   _zz_750;
  wire       [0:0]    _zz_751;
  wire       [0:0]    _zz_752;
  wire       [15:0]   _zz_753;
  wire       [15:0]   _zz_754;
  wire       [0:0]    _zz_755;
  wire       [0:0]    _zz_756;
  wire       [15:0]   _zz_757;
  wire       [15:0]   _zz_758;
  wire       [0:0]    _zz_759;
  wire       [0:0]    _zz_760;
  wire       [15:0]   _zz_761;
  wire       [15:0]   _zz_762;
  wire       [0:0]    _zz_763;
  wire       [0:0]    _zz_764;
  wire       [15:0]   _zz_765;
  wire       [15:0]   _zz_766;
  wire       [0:0]    _zz_767;
  wire       [0:0]    _zz_768;
  wire       [15:0]   _zz_769;
  wire       [15:0]   _zz_770;
  wire       [0:0]    _zz_771;
  wire       [0:0]    _zz_772;
  wire       [15:0]   _zz_773;
  wire       [15:0]   _zz_774;
  wire       [0:0]    _zz_775;
  wire       [0:0]    _zz_776;
  wire       [15:0]   _zz_777;
  wire       [15:0]   _zz_778;
  wire       [0:0]    _zz_779;
  wire       [0:0]    _zz_780;
  wire       [15:0]   _zz_781;
  wire       [15:0]   _zz_782;
  wire       [0:0]    _zz_783;
  wire       [0:0]    _zz_784;
  wire       [15:0]   _zz_785;
  wire       [15:0]   _zz_786;
  wire       [0:0]    _zz_787;
  wire       [0:0]    _zz_788;
  wire       [15:0]   _zz_789;
  wire       [15:0]   _zz_790;
  wire       [0:0]    _zz_791;
  wire       [0:0]    _zz_792;
  wire       [15:0]   _zz_793;
  wire       [15:0]   _zz_794;
  wire       [0:0]    _zz_795;
  wire       [0:0]    _zz_796;
  wire       [15:0]   _zz_797;
  wire       [15:0]   _zz_798;
  wire       [0:0]    _zz_799;
  wire       [0:0]    _zz_800;
  wire       [15:0]   _zz_801;
  wire       [15:0]   _zz_802;
  wire       [0:0]    _zz_803;
  wire       [0:0]    _zz_804;
  wire       [15:0]   _zz_805;
  wire       [15:0]   _zz_806;
  wire       [0:0]    _zz_807;
  wire       [0:0]    _zz_808;
  wire       [15:0]   _zz_809;
  wire       [15:0]   _zz_810;
  wire       [0:0]    _zz_811;
  wire       [0:0]    _zz_812;
  wire       [15:0]   _zz_813;
  wire       [15:0]   _zz_814;
  wire       [0:0]    _zz_815;
  wire       [0:0]    _zz_816;
  wire       [15:0]   _zz_817;
  wire       [15:0]   _zz_818;
  wire       [0:0]    _zz_819;
  wire       [0:0]    _zz_820;
  wire       [15:0]   _zz_821;
  wire       [15:0]   _zz_822;
  wire       [0:0]    _zz_823;
  wire       [0:0]    _zz_824;
  wire       [15:0]   _zz_825;
  wire       [15:0]   _zz_826;
  wire       [0:0]    _zz_827;
  wire       [0:0]    _zz_828;
  wire       [15:0]   _zz_829;
  wire       [15:0]   _zz_830;
  wire       [0:0]    _zz_831;
  wire       [0:0]    _zz_832;
  wire       [15:0]   _zz_833;
  wire       [15:0]   _zz_834;
  wire       [0:0]    _zz_835;
  wire       [0:0]    _zz_836;
  wire       [15:0]   _zz_837;
  wire       [15:0]   _zz_838;
  wire       [0:0]    _zz_839;
  wire       [0:0]    _zz_840;
  wire       [15:0]   _zz_841;
  wire       [15:0]   _zz_842;
  wire       [0:0]    _zz_843;
  wire       [0:0]    _zz_844;
  wire       [15:0]   _zz_845;
  wire       [15:0]   _zz_846;
  wire       [0:0]    _zz_847;
  wire       [0:0]    _zz_848;
  wire       [15:0]   _zz_849;
  wire       [15:0]   _zz_850;
  wire       [0:0]    _zz_851;
  wire       [0:0]    _zz_852;
  wire       [15:0]   _zz_853;
  wire       [15:0]   _zz_854;
  wire       [0:0]    _zz_855;
  wire       [0:0]    _zz_856;
  wire       [15:0]   _zz_857;
  wire       [15:0]   _zz_858;
  wire       [0:0]    _zz_859;
  wire       [0:0]    _zz_860;
  wire       [15:0]   _zz_861;
  wire       [15:0]   _zz_862;
  wire       [0:0]    _zz_863;
  wire       [0:0]    _zz_864;
  wire       [15:0]   _zz_865;
  wire       [15:0]   _zz_866;
  wire       [0:0]    _zz_867;
  wire       [0:0]    _zz_868;
  wire       [15:0]   _zz_869;
  wire       [15:0]   _zz_870;
  wire       [0:0]    _zz_871;
  wire       [0:0]    _zz_872;
  wire       [15:0]   _zz_873;
  wire       [15:0]   _zz_874;
  wire       [0:0]    _zz_875;
  wire       [0:0]    _zz_876;
  wire       [15:0]   _zz_877;
  wire       [15:0]   _zz_878;
  wire       [0:0]    _zz_879;
  wire       [0:0]    _zz_880;
  wire       [15:0]   _zz_881;
  wire       [15:0]   _zz_882;
  wire       [0:0]    _zz_883;
  wire       [0:0]    _zz_884;
  wire       [15:0]   _zz_885;
  wire       [15:0]   _zz_886;
  wire       [0:0]    _zz_887;
  wire       [0:0]    _zz_888;
  wire       [15:0]   _zz_889;
  wire       [15:0]   _zz_890;
  wire       [0:0]    _zz_891;
  wire       [0:0]    _zz_892;
  wire       [15:0]   _zz_893;
  wire       [15:0]   _zz_894;
  wire       [0:0]    _zz_895;
  wire       [0:0]    _zz_896;
  wire       [15:0]   _zz_897;
  wire       [15:0]   _zz_898;
  wire       [0:0]    _zz_899;
  wire       [0:0]    _zz_900;
  wire       [15:0]   _zz_901;
  wire       [15:0]   _zz_902;
  wire       [0:0]    _zz_903;
  wire       [0:0]    _zz_904;
  wire       [15:0]   _zz_905;
  wire       [15:0]   _zz_906;
  wire       [0:0]    _zz_907;
  wire       [0:0]    _zz_908;
  wire       [15:0]   _zz_909;
  wire       [15:0]   _zz_910;
  wire       [0:0]    _zz_911;
  wire       [0:0]    _zz_912;
  wire       [15:0]   _zz_913;
  wire       [15:0]   _zz_914;
  wire       [0:0]    _zz_915;
  wire       [0:0]    _zz_916;
  wire       [15:0]   _zz_917;
  wire       [15:0]   _zz_918;
  wire       [0:0]    _zz_919;
  wire       [0:0]    _zz_920;
  wire       [15:0]   _zz_921;
  wire       [15:0]   _zz_922;
  wire       [0:0]    _zz_923;
  wire       [0:0]    _zz_924;
  wire       [15:0]   _zz_925;
  wire       [15:0]   _zz_926;
  wire       [0:0]    _zz_927;
  wire       [0:0]    _zz_928;
  wire       [15:0]   _zz_929;
  wire       [15:0]   _zz_930;
  wire       [0:0]    _zz_931;
  wire       [0:0]    _zz_932;
  wire       [15:0]   _zz_933;
  wire       [15:0]   _zz_934;
  wire       [0:0]    _zz_935;
  wire       [0:0]    _zz_936;
  wire       [15:0]   _zz_937;
  wire       [15:0]   _zz_938;
  wire       [0:0]    _zz_939;
  wire       [0:0]    _zz_940;
  wire       [15:0]   _zz_941;
  wire       [15:0]   _zz_942;
  wire       [0:0]    _zz_943;
  wire       [0:0]    _zz_944;
  wire       [15:0]   _zz_945;
  wire       [15:0]   _zz_946;
  wire       [0:0]    _zz_947;
  wire       [0:0]    _zz_948;
  wire       [15:0]   _zz_949;
  wire       [15:0]   _zz_950;
  wire       [0:0]    _zz_951;
  wire       [0:0]    _zz_952;
  wire       [15:0]   _zz_953;
  wire       [15:0]   _zz_954;
  wire       [0:0]    _zz_955;
  wire       [0:0]    _zz_956;
  wire       [15:0]   _zz_957;
  wire       [15:0]   _zz_958;
  wire       [0:0]    _zz_959;
  wire       [0:0]    _zz_960;
  wire       [15:0]   _zz_961;
  wire       [15:0]   _zz_962;
  wire       [0:0]    _zz_963;
  wire       [0:0]    _zz_964;
  wire       [15:0]   _zz_965;
  wire       [15:0]   _zz_966;
  wire       [0:0]    _zz_967;
  wire       [0:0]    _zz_968;
  wire       [15:0]   _zz_969;
  wire       [15:0]   _zz_970;
  wire       [0:0]    _zz_971;
  wire       [0:0]    _zz_972;
  wire       [15:0]   _zz_973;
  wire       [15:0]   _zz_974;
  wire       [0:0]    _zz_975;
  wire       [0:0]    _zz_976;
  wire       [15:0]   _zz_977;
  wire       [15:0]   _zz_978;
  wire       [0:0]    _zz_979;
  wire       [0:0]    _zz_980;
  wire       [15:0]   _zz_981;
  wire       [15:0]   _zz_982;
  wire       [0:0]    _zz_983;
  wire       [0:0]    _zz_984;
  wire       [15:0]   _zz_985;
  wire       [15:0]   _zz_986;
  wire       [0:0]    _zz_987;
  wire       [0:0]    _zz_988;
  wire       [15:0]   _zz_989;
  wire       [15:0]   _zz_990;
  wire       [0:0]    _zz_991;
  wire       [0:0]    _zz_992;
  wire       [15:0]   _zz_993;
  wire       [15:0]   _zz_994;
  wire       [0:0]    _zz_995;
  wire       [0:0]    _zz_996;
  wire       [15:0]   _zz_997;
  wire       [15:0]   _zz_998;
  wire       [0:0]    _zz_999;
  wire       [0:0]    _zz_1000;
  wire       [15:0]   _zz_1001;
  wire       [15:0]   _zz_1002;
  wire       [0:0]    _zz_1003;
  wire       [0:0]    _zz_1004;
  wire       [15:0]   _zz_1005;
  wire       [15:0]   _zz_1006;
  wire       [0:0]    _zz_1007;
  wire       [0:0]    _zz_1008;
  wire       [15:0]   _zz_1009;
  wire       [15:0]   _zz_1010;
  wire       [0:0]    _zz_1011;
  wire       [0:0]    _zz_1012;
  wire       [15:0]   _zz_1013;
  wire       [15:0]   _zz_1014;
  wire       [0:0]    _zz_1015;
  wire       [0:0]    _zz_1016;
  wire       [15:0]   _zz_1017;
  wire       [15:0]   _zz_1018;
  wire       [0:0]    _zz_1019;
  wire       [0:0]    _zz_1020;
  wire       [15:0]   _zz_1021;
  wire       [15:0]   _zz_1022;
  wire       [0:0]    _zz_1023;
  wire       [0:0]    _zz_1024;
  wire       [15:0]   _zz_1025;
  wire       [15:0]   _zz_1026;
  wire       [0:0]    _zz_1027;
  wire       [0:0]    _zz_1028;
  wire       [15:0]   _zz_1029;
  wire       [15:0]   _zz_1030;
  wire       [0:0]    _zz_1031;
  wire       [0:0]    _zz_1032;
  wire       [15:0]   _zz_1033;
  wire       [15:0]   _zz_1034;
  wire       [0:0]    _zz_1035;
  wire       [0:0]    _zz_1036;
  wire       [15:0]   _zz_1037;
  wire       [15:0]   _zz_1038;
  wire       [0:0]    _zz_1039;
  wire       [0:0]    _zz_1040;
  wire       [15:0]   _zz_1041;
  wire       [15:0]   _zz_1042;
  wire       [0:0]    _zz_1043;
  wire       [0:0]    _zz_1044;
  wire       [15:0]   _zz_1045;
  wire       [15:0]   _zz_1046;
  wire       [0:0]    _zz_1047;
  wire       [0:0]    _zz_1048;
  wire       [15:0]   _zz_1049;
  wire       [15:0]   _zz_1050;
  wire       [0:0]    _zz_1051;
  wire       [0:0]    _zz_1052;
  wire       [15:0]   _zz_1053;
  wire       [15:0]   _zz_1054;
  wire       [0:0]    _zz_1055;
  wire       [0:0]    _zz_1056;
  wire       [15:0]   _zz_1057;
  wire       [15:0]   _zz_1058;
  wire       [0:0]    _zz_1059;
  wire       [0:0]    _zz_1060;
  wire       [15:0]   _zz_1061;
  wire       [15:0]   _zz_1062;
  wire       [0:0]    _zz_1063;
  wire       [0:0]    _zz_1064;
  wire       [15:0]   _zz_1065;
  wire       [15:0]   _zz_1066;
  wire       [0:0]    _zz_1067;
  wire       [0:0]    _zz_1068;
  wire       [15:0]   _zz_1069;
  wire       [15:0]   _zz_1070;
  wire       [0:0]    _zz_1071;
  wire       [0:0]    _zz_1072;
  wire       [15:0]   _zz_1073;
  wire       [15:0]   _zz_1074;
  wire       [0:0]    _zz_1075;
  wire       [0:0]    _zz_1076;
  wire       [15:0]   _zz_1077;
  wire       [15:0]   _zz_1078;
  wire       [0:0]    _zz_1079;
  wire       [0:0]    _zz_1080;
  wire       [15:0]   _zz_1081;
  wire       [15:0]   _zz_1082;
  wire       [0:0]    _zz_1083;
  wire       [0:0]    _zz_1084;
  wire       [15:0]   _zz_1085;
  wire       [15:0]   _zz_1086;
  wire       [0:0]    _zz_1087;
  wire       [0:0]    _zz_1088;
  wire       [15:0]   _zz_1089;
  wire       [15:0]   _zz_1090;
  wire       [0:0]    _zz_1091;
  wire       [0:0]    _zz_1092;
  wire       [15:0]   _zz_1093;
  wire       [15:0]   _zz_1094;
  wire       [0:0]    _zz_1095;
  wire       [0:0]    _zz_1096;
  wire       [15:0]   _zz_1097;
  wire       [15:0]   _zz_1098;
  wire       [0:0]    _zz_1099;
  wire       [0:0]    _zz_1100;
  wire       [15:0]   _zz_1101;
  wire       [15:0]   _zz_1102;
  wire       [0:0]    _zz_1103;
  wire       [0:0]    _zz_1104;
  wire       [15:0]   _zz_1105;
  wire       [15:0]   _zz_1106;
  wire       [0:0]    _zz_1107;
  wire       [0:0]    _zz_1108;
  wire       [15:0]   _zz_1109;
  wire       [15:0]   _zz_1110;
  wire       [0:0]    _zz_1111;
  wire       [0:0]    _zz_1112;
  wire       [15:0]   _zz_1113;
  wire       [15:0]   _zz_1114;
  wire       [0:0]    _zz_1115;
  wire       [0:0]    _zz_1116;
  wire       [15:0]   _zz_1117;
  wire       [15:0]   _zz_1118;
  wire       [0:0]    _zz_1119;
  wire       [0:0]    _zz_1120;
  wire       [15:0]   _zz_1121;
  wire       [15:0]   _zz_1122;
  wire       [0:0]    _zz_1123;
  wire       [0:0]    _zz_1124;
  wire       [15:0]   _zz_1125;
  wire       [15:0]   _zz_1126;
  wire       [0:0]    _zz_1127;
  wire       [0:0]    _zz_1128;
  wire       [15:0]   _zz_1129;
  wire       [15:0]   _zz_1130;
  wire       [0:0]    _zz_1131;
  wire       [0:0]    _zz_1132;
  wire       [15:0]   _zz_1133;
  wire       [15:0]   _zz_1134;
  wire       [0:0]    _zz_1135;
  wire       [0:0]    _zz_1136;
  wire       [15:0]   _zz_1137;
  wire       [15:0]   _zz_1138;
  wire       [0:0]    _zz_1139;
  wire       [0:0]    _zz_1140;
  wire       [15:0]   _zz_1141;
  wire       [15:0]   _zz_1142;
  wire       [0:0]    _zz_1143;
  wire       [0:0]    _zz_1144;
  wire       [15:0]   _zz_1145;
  wire       [15:0]   _zz_1146;
  wire       [0:0]    _zz_1147;
  wire       [0:0]    _zz_1148;
  wire       [15:0]   _zz_1149;
  wire       [15:0]   _zz_1150;
  wire       [0:0]    _zz_1151;
  wire       [0:0]    _zz_1152;
  wire       [15:0]   _zz_1153;
  wire       [15:0]   _zz_1154;
  wire       [0:0]    _zz_1155;
  wire       [0:0]    _zz_1156;
  wire       [15:0]   _zz_1157;
  wire       [15:0]   _zz_1158;
  wire       [0:0]    _zz_1159;
  wire       [0:0]    _zz_1160;
  wire       [15:0]   _zz_1161;
  wire       [15:0]   _zz_1162;
  wire       [0:0]    _zz_1163;
  wire       [0:0]    _zz_1164;
  wire       [15:0]   _zz_1165;
  wire       [15:0]   _zz_1166;
  wire       [0:0]    _zz_1167;
  wire       [0:0]    _zz_1168;
  wire       [15:0]   _zz_1169;
  wire       [15:0]   _zz_1170;
  wire       [0:0]    _zz_1171;
  wire       [0:0]    _zz_1172;
  wire       [15:0]   _zz_1173;
  wire       [15:0]   _zz_1174;
  wire       [0:0]    _zz_1175;
  wire       [0:0]    _zz_1176;
  wire       [15:0]   _zz_1177;
  wire       [15:0]   _zz_1178;
  wire       [0:0]    _zz_1179;
  wire       [0:0]    _zz_1180;
  wire       [15:0]   _zz_1181;
  wire       [15:0]   _zz_1182;
  wire       [0:0]    _zz_1183;
  wire       [0:0]    _zz_1184;
  wire       [15:0]   _zz_1185;
  wire       [15:0]   _zz_1186;
  wire       [0:0]    _zz_1187;
  wire       [0:0]    _zz_1188;
  wire       [15:0]   _zz_1189;
  wire       [15:0]   _zz_1190;
  wire       [0:0]    _zz_1191;
  wire       [0:0]    _zz_1192;
  wire       [15:0]   _zz_1193;
  wire       [15:0]   _zz_1194;
  wire       [0:0]    _zz_1195;
  wire       [0:0]    _zz_1196;
  wire       [15:0]   _zz_1197;
  wire       [15:0]   _zz_1198;
  wire       [0:0]    _zz_1199;
  wire       [0:0]    _zz_1200;
  wire       [15:0]   _zz_1201;
  wire       [15:0]   _zz_1202;
  wire       [0:0]    _zz_1203;
  wire       [0:0]    _zz_1204;
  wire       [15:0]   _zz_1205;
  wire       [15:0]   _zz_1206;
  wire       [0:0]    _zz_1207;
  wire       [0:0]    _zz_1208;
  wire       [15:0]   _zz_1209;
  wire       [15:0]   _zz_1210;
  wire       [0:0]    _zz_1211;
  wire       [0:0]    _zz_1212;
  wire       [15:0]   _zz_1213;
  wire       [15:0]   _zz_1214;
  wire       [0:0]    _zz_1215;
  wire       [0:0]    _zz_1216;
  wire       [15:0]   _zz_1217;
  wire       [15:0]   _zz_1218;
  wire       [0:0]    _zz_1219;
  wire       [0:0]    _zz_1220;
  wire       [15:0]   _zz_1221;
  wire       [15:0]   _zz_1222;
  wire       [0:0]    _zz_1223;
  wire       [0:0]    _zz_1224;
  wire       [15:0]   _zz_1225;
  wire       [15:0]   _zz_1226;
  wire       [0:0]    _zz_1227;
  wire       [0:0]    _zz_1228;
  wire       [15:0]   _zz_1229;
  wire       [15:0]   _zz_1230;
  wire       [0:0]    _zz_1231;
  wire       [0:0]    _zz_1232;
  wire       [15:0]   _zz_1233;
  wire       [15:0]   _zz_1234;
  wire       [0:0]    _zz_1235;
  wire       [0:0]    _zz_1236;
  wire       [15:0]   _zz_1237;
  wire       [15:0]   _zz_1238;
  wire       [0:0]    _zz_1239;
  wire       [0:0]    _zz_1240;
  wire       [15:0]   _zz_1241;
  wire       [15:0]   _zz_1242;
  wire       [0:0]    _zz_1243;
  wire       [0:0]    _zz_1244;
  wire       [15:0]   _zz_1245;
  wire       [15:0]   _zz_1246;
  wire       [0:0]    _zz_1247;
  wire       [0:0]    _zz_1248;
  wire       [15:0]   _zz_1249;
  wire       [15:0]   _zz_1250;
  wire       [0:0]    _zz_1251;
  wire       [0:0]    _zz_1252;
  wire       [15:0]   _zz_1253;
  wire       [15:0]   _zz_1254;
  wire       [0:0]    _zz_1255;
  wire       [0:0]    _zz_1256;
  wire       [15:0]   _zz_1257;
  wire       [15:0]   _zz_1258;
  wire       [0:0]    _zz_1259;
  wire       [0:0]    _zz_1260;
  wire       [15:0]   _zz_1261;
  wire       [15:0]   _zz_1262;
  wire       [0:0]    _zz_1263;
  wire       [0:0]    _zz_1264;
  wire       [15:0]   _zz_1265;
  wire       [15:0]   _zz_1266;
  wire       [0:0]    _zz_1267;
  wire       [0:0]    _zz_1268;
  wire       [15:0]   _zz_1269;
  wire       [15:0]   _zz_1270;
  wire       [0:0]    _zz_1271;
  wire       [0:0]    _zz_1272;
  wire       [15:0]   _zz_1273;
  wire       [15:0]   _zz_1274;
  wire       [0:0]    _zz_1275;
  wire       [0:0]    _zz_1276;
  wire       [15:0]   _zz_1277;
  wire       [15:0]   _zz_1278;
  wire       [0:0]    _zz_1279;
  wire       [0:0]    _zz_1280;
  wire       [15:0]   _zz_1281;
  wire       [15:0]   _zz_1282;
  wire       [0:0]    _zz_1283;
  wire       [0:0]    _zz_1284;
  wire       [15:0]   _zz_1285;
  wire       [15:0]   _zz_1286;
  wire       [0:0]    _zz_1287;
  wire       [0:0]    _zz_1288;
  wire       [15:0]   _zz_1289;
  wire       [15:0]   _zz_1290;
  wire       [0:0]    _zz_1291;
  wire       [0:0]    _zz_1292;
  wire       [15:0]   _zz_1293;
  wire       [15:0]   _zz_1294;
  wire       [0:0]    _zz_1295;
  wire       [0:0]    _zz_1296;
  wire       [15:0]   _zz_1297;
  wire       [15:0]   _zz_1298;
  wire       [0:0]    _zz_1299;
  wire       [0:0]    _zz_1300;
  wire       [15:0]   _zz_1301;
  wire       [15:0]   _zz_1302;
  wire       [0:0]    _zz_1303;
  wire       [0:0]    _zz_1304;
  wire       [15:0]   _zz_1305;
  wire       [15:0]   _zz_1306;
  wire       [0:0]    _zz_1307;
  wire       [0:0]    _zz_1308;
  wire       [15:0]   _zz_1309;
  wire       [15:0]   _zz_1310;
  wire       [0:0]    _zz_1311;
  wire       [0:0]    _zz_1312;
  wire       [15:0]   _zz_1313;
  wire       [15:0]   _zz_1314;
  wire       [0:0]    _zz_1315;
  wire       [0:0]    _zz_1316;
  wire       [15:0]   _zz_1317;
  wire       [15:0]   _zz_1318;
  wire       [0:0]    _zz_1319;
  wire       [0:0]    _zz_1320;
  wire       [15:0]   _zz_1321;
  wire       [15:0]   _zz_1322;
  wire       [0:0]    _zz_1323;
  wire       [0:0]    _zz_1324;
  wire       [15:0]   _zz_1325;
  wire       [15:0]   _zz_1326;
  wire       [0:0]    _zz_1327;
  wire       [0:0]    _zz_1328;
  wire       [15:0]   _zz_1329;
  wire       [15:0]   _zz_1330;
  wire       [0:0]    _zz_1331;
  wire       [0:0]    _zz_1332;
  wire       [15:0]   _zz_1333;
  wire       [15:0]   _zz_1334;
  wire       [0:0]    _zz_1335;
  wire       [0:0]    _zz_1336;
  wire       [15:0]   _zz_1337;
  wire       [15:0]   _zz_1338;
  wire       [0:0]    _zz_1339;
  wire       [0:0]    _zz_1340;
  wire       [15:0]   _zz_1341;
  wire       [15:0]   _zz_1342;
  wire       [0:0]    _zz_1343;
  wire       [0:0]    _zz_1344;
  wire       [15:0]   _zz_1345;
  wire       [15:0]   _zz_1346;
  wire       [0:0]    _zz_1347;
  wire       [0:0]    _zz_1348;
  wire       [15:0]   _zz_1349;
  wire       [15:0]   _zz_1350;
  wire       [0:0]    _zz_1351;
  wire       [0:0]    _zz_1352;
  wire       [15:0]   _zz_1353;
  wire       [15:0]   _zz_1354;
  wire       [0:0]    _zz_1355;
  wire       [0:0]    _zz_1356;
  wire       [15:0]   _zz_1357;
  wire       [15:0]   _zz_1358;
  wire       [0:0]    _zz_1359;
  wire       [0:0]    _zz_1360;
  wire       [15:0]   _zz_1361;
  wire       [15:0]   _zz_1362;
  wire       [0:0]    _zz_1363;
  wire       [0:0]    _zz_1364;
  wire       [15:0]   _zz_1365;
  wire       [15:0]   _zz_1366;
  wire       [0:0]    _zz_1367;
  wire       [0:0]    _zz_1368;
  wire       [15:0]   _zz_1369;
  wire       [15:0]   _zz_1370;
  wire       [0:0]    _zz_1371;
  wire       [0:0]    _zz_1372;
  wire       [15:0]   _zz_1373;
  wire       [15:0]   _zz_1374;
  wire       [0:0]    _zz_1375;
  wire       [0:0]    _zz_1376;
  wire       [15:0]   _zz_1377;
  wire       [15:0]   _zz_1378;
  wire       [0:0]    _zz_1379;
  wire       [0:0]    _zz_1380;
  wire       [15:0]   _zz_1381;
  wire       [15:0]   _zz_1382;
  wire       [0:0]    _zz_1383;
  wire       [0:0]    _zz_1384;
  wire       [15:0]   _zz_1385;
  wire       [15:0]   _zz_1386;
  wire       [0:0]    _zz_1387;
  wire       [0:0]    _zz_1388;
  wire       [15:0]   _zz_1389;
  wire       [15:0]   _zz_1390;
  wire       [0:0]    _zz_1391;
  wire       [0:0]    _zz_1392;
  wire       [15:0]   _zz_1393;
  wire       [15:0]   _zz_1394;
  wire       [0:0]    _zz_1395;
  wire       [0:0]    _zz_1396;
  wire       [15:0]   _zz_1397;
  wire       [15:0]   _zz_1398;
  wire       [0:0]    _zz_1399;
  wire       [0:0]    _zz_1400;
  wire       [15:0]   _zz_1401;
  wire       [15:0]   _zz_1402;
  wire       [0:0]    _zz_1403;
  wire       [0:0]    _zz_1404;
  wire       [15:0]   _zz_1405;
  wire       [15:0]   _zz_1406;
  wire       [0:0]    _zz_1407;
  wire       [0:0]    _zz_1408;
  wire       [15:0]   _zz_1409;
  wire       [15:0]   _zz_1410;
  wire       [0:0]    _zz_1411;
  wire       [0:0]    _zz_1412;
  wire       [15:0]   _zz_1413;
  wire       [15:0]   _zz_1414;
  wire       [0:0]    _zz_1415;
  wire       [0:0]    _zz_1416;
  wire       [15:0]   _zz_1417;
  wire       [15:0]   _zz_1418;
  wire       [0:0]    _zz_1419;
  wire       [0:0]    _zz_1420;
  wire       [15:0]   _zz_1421;
  wire       [15:0]   _zz_1422;
  wire       [0:0]    _zz_1423;
  wire       [0:0]    _zz_1424;
  wire       [15:0]   _zz_1425;
  wire       [15:0]   _zz_1426;
  wire       [0:0]    _zz_1427;
  wire       [0:0]    _zz_1428;
  wire       [15:0]   _zz_1429;
  wire       [15:0]   _zz_1430;
  wire       [0:0]    _zz_1431;
  wire       [0:0]    _zz_1432;
  wire       [15:0]   _zz_1433;
  wire       [15:0]   _zz_1434;
  wire       [0:0]    _zz_1435;
  wire       [0:0]    _zz_1436;
  wire       [15:0]   _zz_1437;
  wire       [15:0]   _zz_1438;
  wire       [0:0]    _zz_1439;
  wire       [0:0]    _zz_1440;
  wire       [15:0]   _zz_1441;
  wire       [15:0]   _zz_1442;
  wire       [0:0]    _zz_1443;
  wire       [0:0]    _zz_1444;
  wire       [15:0]   _zz_1445;
  wire       [15:0]   _zz_1446;
  wire       [0:0]    _zz_1447;
  wire       [0:0]    _zz_1448;
  wire       [15:0]   _zz_1449;
  wire       [15:0]   _zz_1450;
  wire       [0:0]    _zz_1451;
  wire       [0:0]    _zz_1452;
  wire       [15:0]   _zz_1453;
  wire       [15:0]   _zz_1454;
  wire       [0:0]    _zz_1455;
  wire       [0:0]    _zz_1456;
  wire       [15:0]   _zz_1457;
  wire       [15:0]   _zz_1458;
  wire       [0:0]    _zz_1459;
  wire       [0:0]    _zz_1460;
  wire       [15:0]   _zz_1461;
  wire       [15:0]   _zz_1462;
  wire       [0:0]    _zz_1463;
  wire       [0:0]    _zz_1464;
  wire       [15:0]   _zz_1465;
  wire       [15:0]   _zz_1466;
  wire       [0:0]    _zz_1467;
  wire       [0:0]    _zz_1468;
  wire       [15:0]   _zz_1469;
  wire       [15:0]   _zz_1470;
  wire       [0:0]    _zz_1471;
  wire       [0:0]    _zz_1472;
  wire       [15:0]   _zz_1473;
  wire       [15:0]   _zz_1474;
  wire       [0:0]    _zz_1475;
  wire       [0:0]    _zz_1476;
  wire       [15:0]   _zz_1477;
  wire       [15:0]   _zz_1478;
  wire       [0:0]    _zz_1479;
  wire       [0:0]    _zz_1480;
  wire       [15:0]   _zz_1481;
  wire       [15:0]   _zz_1482;
  wire       [0:0]    _zz_1483;
  wire       [0:0]    _zz_1484;
  wire       [15:0]   _zz_1485;
  wire       [15:0]   _zz_1486;
  wire       [0:0]    _zz_1487;
  wire       [0:0]    _zz_1488;
  wire       [15:0]   _zz_1489;
  wire       [15:0]   _zz_1490;
  wire       [0:0]    _zz_1491;
  wire       [0:0]    _zz_1492;
  wire       [15:0]   _zz_1493;
  wire       [15:0]   _zz_1494;
  wire       [0:0]    _zz_1495;
  wire       [0:0]    _zz_1496;
  wire       [15:0]   _zz_1497;
  wire       [15:0]   _zz_1498;
  wire       [0:0]    _zz_1499;
  wire       [0:0]    _zz_1500;
  wire       [15:0]   _zz_1501;
  wire       [15:0]   _zz_1502;
  wire       [0:0]    _zz_1503;
  wire       [0:0]    _zz_1504;
  wire       [15:0]   _zz_1505;
  wire       [15:0]   _zz_1506;
  wire       [0:0]    _zz_1507;
  wire       [0:0]    _zz_1508;
  wire       [15:0]   _zz_1509;
  wire       [15:0]   _zz_1510;
  wire       [0:0]    _zz_1511;
  wire       [0:0]    _zz_1512;
  wire       [15:0]   _zz_1513;
  wire       [15:0]   _zz_1514;
  wire       [0:0]    _zz_1515;
  wire       [0:0]    _zz_1516;
  wire       [15:0]   _zz_1517;
  wire       [15:0]   _zz_1518;
  wire       [0:0]    _zz_1519;
  wire       [0:0]    _zz_1520;
  wire       [15:0]   _zz_1521;
  wire       [15:0]   _zz_1522;
  wire       [0:0]    _zz_1523;
  wire       [0:0]    _zz_1524;
  wire       [15:0]   _zz_1525;
  wire       [15:0]   _zz_1526;
  wire       [0:0]    _zz_1527;
  wire       [0:0]    _zz_1528;
  wire       [15:0]   _zz_1529;
  wire       [15:0]   _zz_1530;
  wire       [0:0]    _zz_1531;
  wire       [0:0]    _zz_1532;
  wire       [15:0]   _zz_1533;
  wire       [15:0]   _zz_1534;
  wire       [0:0]    _zz_1535;
  wire       [0:0]    _zz_1536;
  wire       [15:0]   _zz_1537;
  wire       [15:0]   _zz_1538;
  wire       [0:0]    _zz_1539;
  wire       [0:0]    _zz_1540;
  wire       [15:0]   _zz_1541;
  wire       [15:0]   _zz_1542;
  wire       [0:0]    _zz_1543;
  wire       [0:0]    _zz_1544;
  wire       [15:0]   _zz_1545;
  wire       [15:0]   _zz_1546;
  wire       [0:0]    _zz_1547;
  wire       [0:0]    _zz_1548;
  wire       [15:0]   _zz_1549;
  wire       [15:0]   _zz_1550;
  wire       [0:0]    _zz_1551;
  wire       [0:0]    _zz_1552;
  wire       [15:0]   _zz_1553;
  wire       [15:0]   _zz_1554;
  wire       [0:0]    _zz_1555;
  wire       [0:0]    _zz_1556;
  wire       [15:0]   _zz_1557;
  wire       [15:0]   _zz_1558;
  wire       [0:0]    _zz_1559;
  wire       [0:0]    _zz_1560;
  wire       [15:0]   _zz_1561;
  wire       [15:0]   _zz_1562;
  wire       [0:0]    _zz_1563;
  wire       [0:0]    _zz_1564;
  wire       [15:0]   _zz_1565;
  wire       [15:0]   _zz_1566;
  wire       [0:0]    _zz_1567;
  wire       [0:0]    _zz_1568;
  wire       [15:0]   _zz_1569;
  wire       [15:0]   _zz_1570;
  wire       [0:0]    _zz_1571;
  wire       [0:0]    _zz_1572;
  wire       [15:0]   _zz_1573;
  wire       [15:0]   _zz_1574;
  wire       [0:0]    _zz_1575;
  wire       [0:0]    _zz_1576;
  wire       [15:0]   _zz_1577;
  wire       [15:0]   _zz_1578;
  wire       [0:0]    _zz_1579;
  wire       [0:0]    _zz_1580;
  wire       [15:0]   _zz_1581;
  wire       [15:0]   _zz_1582;
  wire       [0:0]    _zz_1583;
  wire       [0:0]    _zz_1584;
  wire       [15:0]   _zz_1585;
  wire       [15:0]   _zz_1586;
  wire       [0:0]    _zz_1587;
  wire       [0:0]    _zz_1588;
  wire       [15:0]   _zz_1589;
  wire       [15:0]   _zz_1590;
  wire       [0:0]    _zz_1591;
  wire       [0:0]    _zz_1592;
  wire       [15:0]   _zz_1593;
  wire       [15:0]   _zz_1594;
  wire       [0:0]    _zz_1595;
  wire       [0:0]    _zz_1596;
  wire       [15:0]   _zz_1597;
  wire       [15:0]   _zz_1598;
  wire       [0:0]    _zz_1599;
  wire       [0:0]    _zz_1600;
  wire       [15:0]   _zz_1601;
  wire       [15:0]   _zz_1602;
  wire       [0:0]    _zz_1603;
  wire       [0:0]    _zz_1604;
  wire       [15:0]   _zz_1605;
  wire       [15:0]   _zz_1606;
  wire       [0:0]    _zz_1607;
  wire       [0:0]    _zz_1608;
  wire       [15:0]   _zz_1609;
  wire       [15:0]   _zz_1610;
  wire       [0:0]    _zz_1611;
  wire       [0:0]    _zz_1612;
  wire       [15:0]   _zz_1613;
  wire       [15:0]   _zz_1614;
  wire       [0:0]    _zz_1615;
  wire       [0:0]    _zz_1616;
  wire       [15:0]   _zz_1617;
  wire       [15:0]   _zz_1618;
  wire       [0:0]    _zz_1619;
  wire       [0:0]    _zz_1620;
  wire       [15:0]   _zz_1621;
  wire       [15:0]   _zz_1622;
  wire       [0:0]    _zz_1623;
  wire       [0:0]    _zz_1624;
  wire       [15:0]   _zz_1625;
  wire       [15:0]   _zz_1626;
  wire       [0:0]    _zz_1627;
  wire       [0:0]    _zz_1628;
  wire       [15:0]   _zz_1629;
  wire       [15:0]   _zz_1630;
  wire       [0:0]    _zz_1631;
  wire       [0:0]    _zz_1632;
  wire       [15:0]   _zz_1633;
  wire       [15:0]   _zz_1634;
  wire       [0:0]    _zz_1635;
  wire       [0:0]    _zz_1636;
  wire       [15:0]   _zz_1637;
  wire       [15:0]   _zz_1638;
  wire       [0:0]    _zz_1639;
  wire       [0:0]    _zz_1640;
  wire       [15:0]   _zz_1641;
  wire       [15:0]   _zz_1642;
  wire       [0:0]    _zz_1643;
  wire       [0:0]    _zz_1644;
  wire       [15:0]   _zz_1645;
  wire       [15:0]   _zz_1646;
  wire       [0:0]    _zz_1647;
  wire       [0:0]    _zz_1648;
  wire       [15:0]   _zz_1649;
  wire       [15:0]   _zz_1650;
  wire       [0:0]    _zz_1651;
  wire       [0:0]    _zz_1652;
  wire       [15:0]   _zz_1653;
  wire       [15:0]   _zz_1654;
  wire       [0:0]    _zz_1655;
  wire       [0:0]    _zz_1656;
  wire       [15:0]   _zz_1657;
  wire       [15:0]   _zz_1658;
  wire       [0:0]    _zz_1659;
  wire       [0:0]    _zz_1660;
  wire       [15:0]   _zz_1661;
  wire       [15:0]   _zz_1662;
  wire       [0:0]    _zz_1663;
  wire       [0:0]    _zz_1664;
  wire       [15:0]   _zz_1665;
  wire       [15:0]   _zz_1666;
  wire       [0:0]    _zz_1667;
  wire       [0:0]    _zz_1668;
  wire       [15:0]   _zz_1669;
  wire       [15:0]   _zz_1670;
  wire       [0:0]    _zz_1671;
  wire       [0:0]    _zz_1672;
  wire       [15:0]   _zz_1673;
  wire       [15:0]   _zz_1674;
  wire       [0:0]    _zz_1675;
  wire       [0:0]    _zz_1676;
  wire       [15:0]   _zz_1677;
  wire       [15:0]   _zz_1678;
  wire       [0:0]    _zz_1679;
  wire       [0:0]    _zz_1680;
  wire       [15:0]   _zz_1681;
  wire       [15:0]   _zz_1682;
  wire       [0:0]    _zz_1683;
  wire       [0:0]    _zz_1684;
  wire       [15:0]   _zz_1685;
  wire       [15:0]   _zz_1686;
  wire       [0:0]    _zz_1687;
  wire       [0:0]    _zz_1688;
  wire       [15:0]   _zz_1689;
  wire       [15:0]   _zz_1690;
  wire       [0:0]    _zz_1691;
  wire       [0:0]    _zz_1692;
  wire       [15:0]   _zz_1693;
  wire       [15:0]   _zz_1694;
  wire       [0:0]    _zz_1695;
  wire       [0:0]    _zz_1696;
  wire       [15:0]   _zz_1697;
  wire       [15:0]   _zz_1698;
  wire       [0:0]    _zz_1699;
  wire       [0:0]    _zz_1700;
  wire       [15:0]   _zz_1701;
  wire       [15:0]   _zz_1702;
  wire       [0:0]    _zz_1703;
  wire       [0:0]    _zz_1704;
  wire       [15:0]   _zz_1705;
  wire       [15:0]   _zz_1706;
  wire       [0:0]    _zz_1707;
  wire       [0:0]    _zz_1708;
  wire       [15:0]   _zz_1709;
  wire       [15:0]   _zz_1710;
  wire       [0:0]    _zz_1711;
  wire       [0:0]    _zz_1712;
  wire       [15:0]   _zz_1713;
  wire       [15:0]   _zz_1714;
  wire       [0:0]    _zz_1715;
  wire       [0:0]    _zz_1716;
  wire       [15:0]   _zz_1717;
  wire       [15:0]   _zz_1718;
  wire       [0:0]    _zz_1719;
  wire       [0:0]    _zz_1720;
  wire       [15:0]   _zz_1721;
  wire       [15:0]   _zz_1722;
  wire       [0:0]    _zz_1723;
  wire       [0:0]    _zz_1724;
  wire       [15:0]   _zz_1725;
  wire       [15:0]   _zz_1726;
  wire       [0:0]    _zz_1727;
  wire       [0:0]    _zz_1728;
  wire       [15:0]   _zz_1729;
  wire       [15:0]   _zz_1730;
  wire       [0:0]    _zz_1731;
  wire       [0:0]    _zz_1732;
  wire       [15:0]   _zz_1733;
  wire       [15:0]   _zz_1734;
  wire       [0:0]    _zz_1735;
  wire       [0:0]    _zz_1736;
  wire       [15:0]   _zz_1737;
  wire       [15:0]   _zz_1738;
  wire       [0:0]    _zz_1739;
  wire       [0:0]    _zz_1740;
  wire       [15:0]   _zz_1741;
  wire       [15:0]   _zz_1742;
  wire       [0:0]    _zz_1743;
  wire       [0:0]    _zz_1744;
  wire       [15:0]   _zz_1745;
  wire       [15:0]   _zz_1746;
  wire       [0:0]    _zz_1747;
  wire       [0:0]    _zz_1748;
  wire       [15:0]   _zz_1749;
  wire       [15:0]   _zz_1750;
  wire       [0:0]    _zz_1751;
  wire       [0:0]    _zz_1752;
  wire       [15:0]   _zz_1753;
  wire       [15:0]   _zz_1754;
  wire       [0:0]    _zz_1755;
  wire       [0:0]    _zz_1756;
  wire       [15:0]   _zz_1757;
  wire       [15:0]   _zz_1758;
  wire       [0:0]    _zz_1759;
  wire       [0:0]    _zz_1760;
  wire       [15:0]   _zz_1761;
  wire       [15:0]   _zz_1762;
  wire       [0:0]    _zz_1763;
  wire       [0:0]    _zz_1764;
  wire       [15:0]   _zz_1765;
  wire       [15:0]   _zz_1766;
  wire       [0:0]    _zz_1767;
  wire       [0:0]    _zz_1768;
  wire       [15:0]   _zz_1769;
  wire       [15:0]   _zz_1770;
  wire       [0:0]    _zz_1771;
  wire       [0:0]    _zz_1772;
  wire       [15:0]   _zz_1773;
  wire       [15:0]   _zz_1774;
  wire       [0:0]    _zz_1775;
  wire       [0:0]    _zz_1776;
  wire       [15:0]   _zz_1777;
  wire       [15:0]   _zz_1778;
  wire       [0:0]    _zz_1779;
  wire       [0:0]    _zz_1780;
  wire       [15:0]   _zz_1781;
  wire       [15:0]   _zz_1782;
  wire       [0:0]    _zz_1783;
  wire       [0:0]    _zz_1784;
  wire       [15:0]   _zz_1785;
  wire       [15:0]   _zz_1786;
  wire       [0:0]    _zz_1787;
  wire       [0:0]    _zz_1788;
  wire       [15:0]   _zz_1789;
  wire       [15:0]   _zz_1790;
  wire       [0:0]    _zz_1791;
  wire       [0:0]    _zz_1792;
  reg                 current_level_cnt_willOverflow_regNext;

  assign _zz_2689 = current_level_cnt_willIncrement;
  assign _zz_2690 = {2'd0, _zz_2689};
  assign _zz_2691 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_1_real));
  assign _zz_2692 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_1_imag));
  assign _zz_2693 = fixTo_dout;
  assign _zz_2694 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_1_imag));
  assign _zz_2695 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_1_real));
  assign _zz_2696 = fixTo_1_dout;
  assign _zz_2697 = _zz_2698;
  assign _zz_2698 = ($signed(_zz_2699) >>> _zz_3);
  assign _zz_2699 = _zz_2700;
  assign _zz_2700 = ($signed(data_mid_0_real) - $signed(_zz_1));
  assign _zz_2701 = _zz_2702;
  assign _zz_2702 = ($signed(_zz_2703) >>> _zz_3);
  assign _zz_2703 = _zz_2704;
  assign _zz_2704 = ($signed(data_mid_0_imag) - $signed(_zz_2));
  assign _zz_2705 = _zz_2706;
  assign _zz_2706 = ($signed(_zz_2707) >>> _zz_4);
  assign _zz_2707 = _zz_2708;
  assign _zz_2708 = ($signed(data_mid_0_real) + $signed(_zz_1));
  assign _zz_2709 = _zz_2710;
  assign _zz_2710 = ($signed(_zz_2711) >>> _zz_4);
  assign _zz_2711 = _zz_2712;
  assign _zz_2712 = ($signed(data_mid_0_imag) + $signed(_zz_2));
  assign _zz_2713 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_3_real));
  assign _zz_2714 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_3_imag));
  assign _zz_2715 = fixTo_2_dout;
  assign _zz_2716 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_3_imag));
  assign _zz_2717 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_3_real));
  assign _zz_2718 = fixTo_3_dout;
  assign _zz_2719 = _zz_2720;
  assign _zz_2720 = ($signed(_zz_2721) >>> _zz_7);
  assign _zz_2721 = _zz_2722;
  assign _zz_2722 = ($signed(data_mid_2_real) - $signed(_zz_5));
  assign _zz_2723 = _zz_2724;
  assign _zz_2724 = ($signed(_zz_2725) >>> _zz_7);
  assign _zz_2725 = _zz_2726;
  assign _zz_2726 = ($signed(data_mid_2_imag) - $signed(_zz_6));
  assign _zz_2727 = _zz_2728;
  assign _zz_2728 = ($signed(_zz_2729) >>> _zz_8);
  assign _zz_2729 = _zz_2730;
  assign _zz_2730 = ($signed(data_mid_2_real) + $signed(_zz_5));
  assign _zz_2731 = _zz_2732;
  assign _zz_2732 = ($signed(_zz_2733) >>> _zz_8);
  assign _zz_2733 = _zz_2734;
  assign _zz_2734 = ($signed(data_mid_2_imag) + $signed(_zz_6));
  assign _zz_2735 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_5_real));
  assign _zz_2736 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_5_imag));
  assign _zz_2737 = fixTo_4_dout;
  assign _zz_2738 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_5_imag));
  assign _zz_2739 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_5_real));
  assign _zz_2740 = fixTo_5_dout;
  assign _zz_2741 = _zz_2742;
  assign _zz_2742 = ($signed(_zz_2743) >>> _zz_11);
  assign _zz_2743 = _zz_2744;
  assign _zz_2744 = ($signed(data_mid_4_real) - $signed(_zz_9));
  assign _zz_2745 = _zz_2746;
  assign _zz_2746 = ($signed(_zz_2747) >>> _zz_11);
  assign _zz_2747 = _zz_2748;
  assign _zz_2748 = ($signed(data_mid_4_imag) - $signed(_zz_10));
  assign _zz_2749 = _zz_2750;
  assign _zz_2750 = ($signed(_zz_2751) >>> _zz_12);
  assign _zz_2751 = _zz_2752;
  assign _zz_2752 = ($signed(data_mid_4_real) + $signed(_zz_9));
  assign _zz_2753 = _zz_2754;
  assign _zz_2754 = ($signed(_zz_2755) >>> _zz_12);
  assign _zz_2755 = _zz_2756;
  assign _zz_2756 = ($signed(data_mid_4_imag) + $signed(_zz_10));
  assign _zz_2757 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_7_real));
  assign _zz_2758 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_7_imag));
  assign _zz_2759 = fixTo_6_dout;
  assign _zz_2760 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_7_imag));
  assign _zz_2761 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_7_real));
  assign _zz_2762 = fixTo_7_dout;
  assign _zz_2763 = _zz_2764;
  assign _zz_2764 = ($signed(_zz_2765) >>> _zz_15);
  assign _zz_2765 = _zz_2766;
  assign _zz_2766 = ($signed(data_mid_6_real) - $signed(_zz_13));
  assign _zz_2767 = _zz_2768;
  assign _zz_2768 = ($signed(_zz_2769) >>> _zz_15);
  assign _zz_2769 = _zz_2770;
  assign _zz_2770 = ($signed(data_mid_6_imag) - $signed(_zz_14));
  assign _zz_2771 = _zz_2772;
  assign _zz_2772 = ($signed(_zz_2773) >>> _zz_16);
  assign _zz_2773 = _zz_2774;
  assign _zz_2774 = ($signed(data_mid_6_real) + $signed(_zz_13));
  assign _zz_2775 = _zz_2776;
  assign _zz_2776 = ($signed(_zz_2777) >>> _zz_16);
  assign _zz_2777 = _zz_2778;
  assign _zz_2778 = ($signed(data_mid_6_imag) + $signed(_zz_14));
  assign _zz_2779 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_9_real));
  assign _zz_2780 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_9_imag));
  assign _zz_2781 = fixTo_8_dout;
  assign _zz_2782 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_9_imag));
  assign _zz_2783 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_9_real));
  assign _zz_2784 = fixTo_9_dout;
  assign _zz_2785 = _zz_2786;
  assign _zz_2786 = ($signed(_zz_2787) >>> _zz_19);
  assign _zz_2787 = _zz_2788;
  assign _zz_2788 = ($signed(data_mid_8_real) - $signed(_zz_17));
  assign _zz_2789 = _zz_2790;
  assign _zz_2790 = ($signed(_zz_2791) >>> _zz_19);
  assign _zz_2791 = _zz_2792;
  assign _zz_2792 = ($signed(data_mid_8_imag) - $signed(_zz_18));
  assign _zz_2793 = _zz_2794;
  assign _zz_2794 = ($signed(_zz_2795) >>> _zz_20);
  assign _zz_2795 = _zz_2796;
  assign _zz_2796 = ($signed(data_mid_8_real) + $signed(_zz_17));
  assign _zz_2797 = _zz_2798;
  assign _zz_2798 = ($signed(_zz_2799) >>> _zz_20);
  assign _zz_2799 = _zz_2800;
  assign _zz_2800 = ($signed(data_mid_8_imag) + $signed(_zz_18));
  assign _zz_2801 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_11_real));
  assign _zz_2802 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_11_imag));
  assign _zz_2803 = fixTo_10_dout;
  assign _zz_2804 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_11_imag));
  assign _zz_2805 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_11_real));
  assign _zz_2806 = fixTo_11_dout;
  assign _zz_2807 = _zz_2808;
  assign _zz_2808 = ($signed(_zz_2809) >>> _zz_23);
  assign _zz_2809 = _zz_2810;
  assign _zz_2810 = ($signed(data_mid_10_real) - $signed(_zz_21));
  assign _zz_2811 = _zz_2812;
  assign _zz_2812 = ($signed(_zz_2813) >>> _zz_23);
  assign _zz_2813 = _zz_2814;
  assign _zz_2814 = ($signed(data_mid_10_imag) - $signed(_zz_22));
  assign _zz_2815 = _zz_2816;
  assign _zz_2816 = ($signed(_zz_2817) >>> _zz_24);
  assign _zz_2817 = _zz_2818;
  assign _zz_2818 = ($signed(data_mid_10_real) + $signed(_zz_21));
  assign _zz_2819 = _zz_2820;
  assign _zz_2820 = ($signed(_zz_2821) >>> _zz_24);
  assign _zz_2821 = _zz_2822;
  assign _zz_2822 = ($signed(data_mid_10_imag) + $signed(_zz_22));
  assign _zz_2823 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_13_real));
  assign _zz_2824 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_13_imag));
  assign _zz_2825 = fixTo_12_dout;
  assign _zz_2826 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_13_imag));
  assign _zz_2827 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_13_real));
  assign _zz_2828 = fixTo_13_dout;
  assign _zz_2829 = _zz_2830;
  assign _zz_2830 = ($signed(_zz_2831) >>> _zz_27);
  assign _zz_2831 = _zz_2832;
  assign _zz_2832 = ($signed(data_mid_12_real) - $signed(_zz_25));
  assign _zz_2833 = _zz_2834;
  assign _zz_2834 = ($signed(_zz_2835) >>> _zz_27);
  assign _zz_2835 = _zz_2836;
  assign _zz_2836 = ($signed(data_mid_12_imag) - $signed(_zz_26));
  assign _zz_2837 = _zz_2838;
  assign _zz_2838 = ($signed(_zz_2839) >>> _zz_28);
  assign _zz_2839 = _zz_2840;
  assign _zz_2840 = ($signed(data_mid_12_real) + $signed(_zz_25));
  assign _zz_2841 = _zz_2842;
  assign _zz_2842 = ($signed(_zz_2843) >>> _zz_28);
  assign _zz_2843 = _zz_2844;
  assign _zz_2844 = ($signed(data_mid_12_imag) + $signed(_zz_26));
  assign _zz_2845 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_15_real));
  assign _zz_2846 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_15_imag));
  assign _zz_2847 = fixTo_14_dout;
  assign _zz_2848 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_15_imag));
  assign _zz_2849 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_15_real));
  assign _zz_2850 = fixTo_15_dout;
  assign _zz_2851 = _zz_2852;
  assign _zz_2852 = ($signed(_zz_2853) >>> _zz_31);
  assign _zz_2853 = _zz_2854;
  assign _zz_2854 = ($signed(data_mid_14_real) - $signed(_zz_29));
  assign _zz_2855 = _zz_2856;
  assign _zz_2856 = ($signed(_zz_2857) >>> _zz_31);
  assign _zz_2857 = _zz_2858;
  assign _zz_2858 = ($signed(data_mid_14_imag) - $signed(_zz_30));
  assign _zz_2859 = _zz_2860;
  assign _zz_2860 = ($signed(_zz_2861) >>> _zz_32);
  assign _zz_2861 = _zz_2862;
  assign _zz_2862 = ($signed(data_mid_14_real) + $signed(_zz_29));
  assign _zz_2863 = _zz_2864;
  assign _zz_2864 = ($signed(_zz_2865) >>> _zz_32);
  assign _zz_2865 = _zz_2866;
  assign _zz_2866 = ($signed(data_mid_14_imag) + $signed(_zz_30));
  assign _zz_2867 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_17_real));
  assign _zz_2868 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_17_imag));
  assign _zz_2869 = fixTo_16_dout;
  assign _zz_2870 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_17_imag));
  assign _zz_2871 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_17_real));
  assign _zz_2872 = fixTo_17_dout;
  assign _zz_2873 = _zz_2874;
  assign _zz_2874 = ($signed(_zz_2875) >>> _zz_35);
  assign _zz_2875 = _zz_2876;
  assign _zz_2876 = ($signed(data_mid_16_real) - $signed(_zz_33));
  assign _zz_2877 = _zz_2878;
  assign _zz_2878 = ($signed(_zz_2879) >>> _zz_35);
  assign _zz_2879 = _zz_2880;
  assign _zz_2880 = ($signed(data_mid_16_imag) - $signed(_zz_34));
  assign _zz_2881 = _zz_2882;
  assign _zz_2882 = ($signed(_zz_2883) >>> _zz_36);
  assign _zz_2883 = _zz_2884;
  assign _zz_2884 = ($signed(data_mid_16_real) + $signed(_zz_33));
  assign _zz_2885 = _zz_2886;
  assign _zz_2886 = ($signed(_zz_2887) >>> _zz_36);
  assign _zz_2887 = _zz_2888;
  assign _zz_2888 = ($signed(data_mid_16_imag) + $signed(_zz_34));
  assign _zz_2889 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_19_real));
  assign _zz_2890 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_19_imag));
  assign _zz_2891 = fixTo_18_dout;
  assign _zz_2892 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_19_imag));
  assign _zz_2893 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_19_real));
  assign _zz_2894 = fixTo_19_dout;
  assign _zz_2895 = _zz_2896;
  assign _zz_2896 = ($signed(_zz_2897) >>> _zz_39);
  assign _zz_2897 = _zz_2898;
  assign _zz_2898 = ($signed(data_mid_18_real) - $signed(_zz_37));
  assign _zz_2899 = _zz_2900;
  assign _zz_2900 = ($signed(_zz_2901) >>> _zz_39);
  assign _zz_2901 = _zz_2902;
  assign _zz_2902 = ($signed(data_mid_18_imag) - $signed(_zz_38));
  assign _zz_2903 = _zz_2904;
  assign _zz_2904 = ($signed(_zz_2905) >>> _zz_40);
  assign _zz_2905 = _zz_2906;
  assign _zz_2906 = ($signed(data_mid_18_real) + $signed(_zz_37));
  assign _zz_2907 = _zz_2908;
  assign _zz_2908 = ($signed(_zz_2909) >>> _zz_40);
  assign _zz_2909 = _zz_2910;
  assign _zz_2910 = ($signed(data_mid_18_imag) + $signed(_zz_38));
  assign _zz_2911 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_21_real));
  assign _zz_2912 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_21_imag));
  assign _zz_2913 = fixTo_20_dout;
  assign _zz_2914 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_21_imag));
  assign _zz_2915 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_21_real));
  assign _zz_2916 = fixTo_21_dout;
  assign _zz_2917 = _zz_2918;
  assign _zz_2918 = ($signed(_zz_2919) >>> _zz_43);
  assign _zz_2919 = _zz_2920;
  assign _zz_2920 = ($signed(data_mid_20_real) - $signed(_zz_41));
  assign _zz_2921 = _zz_2922;
  assign _zz_2922 = ($signed(_zz_2923) >>> _zz_43);
  assign _zz_2923 = _zz_2924;
  assign _zz_2924 = ($signed(data_mid_20_imag) - $signed(_zz_42));
  assign _zz_2925 = _zz_2926;
  assign _zz_2926 = ($signed(_zz_2927) >>> _zz_44);
  assign _zz_2927 = _zz_2928;
  assign _zz_2928 = ($signed(data_mid_20_real) + $signed(_zz_41));
  assign _zz_2929 = _zz_2930;
  assign _zz_2930 = ($signed(_zz_2931) >>> _zz_44);
  assign _zz_2931 = _zz_2932;
  assign _zz_2932 = ($signed(data_mid_20_imag) + $signed(_zz_42));
  assign _zz_2933 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_23_real));
  assign _zz_2934 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_23_imag));
  assign _zz_2935 = fixTo_22_dout;
  assign _zz_2936 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_23_imag));
  assign _zz_2937 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_23_real));
  assign _zz_2938 = fixTo_23_dout;
  assign _zz_2939 = _zz_2940;
  assign _zz_2940 = ($signed(_zz_2941) >>> _zz_47);
  assign _zz_2941 = _zz_2942;
  assign _zz_2942 = ($signed(data_mid_22_real) - $signed(_zz_45));
  assign _zz_2943 = _zz_2944;
  assign _zz_2944 = ($signed(_zz_2945) >>> _zz_47);
  assign _zz_2945 = _zz_2946;
  assign _zz_2946 = ($signed(data_mid_22_imag) - $signed(_zz_46));
  assign _zz_2947 = _zz_2948;
  assign _zz_2948 = ($signed(_zz_2949) >>> _zz_48);
  assign _zz_2949 = _zz_2950;
  assign _zz_2950 = ($signed(data_mid_22_real) + $signed(_zz_45));
  assign _zz_2951 = _zz_2952;
  assign _zz_2952 = ($signed(_zz_2953) >>> _zz_48);
  assign _zz_2953 = _zz_2954;
  assign _zz_2954 = ($signed(data_mid_22_imag) + $signed(_zz_46));
  assign _zz_2955 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_25_real));
  assign _zz_2956 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_25_imag));
  assign _zz_2957 = fixTo_24_dout;
  assign _zz_2958 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_25_imag));
  assign _zz_2959 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_25_real));
  assign _zz_2960 = fixTo_25_dout;
  assign _zz_2961 = _zz_2962;
  assign _zz_2962 = ($signed(_zz_2963) >>> _zz_51);
  assign _zz_2963 = _zz_2964;
  assign _zz_2964 = ($signed(data_mid_24_real) - $signed(_zz_49));
  assign _zz_2965 = _zz_2966;
  assign _zz_2966 = ($signed(_zz_2967) >>> _zz_51);
  assign _zz_2967 = _zz_2968;
  assign _zz_2968 = ($signed(data_mid_24_imag) - $signed(_zz_50));
  assign _zz_2969 = _zz_2970;
  assign _zz_2970 = ($signed(_zz_2971) >>> _zz_52);
  assign _zz_2971 = _zz_2972;
  assign _zz_2972 = ($signed(data_mid_24_real) + $signed(_zz_49));
  assign _zz_2973 = _zz_2974;
  assign _zz_2974 = ($signed(_zz_2975) >>> _zz_52);
  assign _zz_2975 = _zz_2976;
  assign _zz_2976 = ($signed(data_mid_24_imag) + $signed(_zz_50));
  assign _zz_2977 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_27_real));
  assign _zz_2978 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_27_imag));
  assign _zz_2979 = fixTo_26_dout;
  assign _zz_2980 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_27_imag));
  assign _zz_2981 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_27_real));
  assign _zz_2982 = fixTo_27_dout;
  assign _zz_2983 = _zz_2984;
  assign _zz_2984 = ($signed(_zz_2985) >>> _zz_55);
  assign _zz_2985 = _zz_2986;
  assign _zz_2986 = ($signed(data_mid_26_real) - $signed(_zz_53));
  assign _zz_2987 = _zz_2988;
  assign _zz_2988 = ($signed(_zz_2989) >>> _zz_55);
  assign _zz_2989 = _zz_2990;
  assign _zz_2990 = ($signed(data_mid_26_imag) - $signed(_zz_54));
  assign _zz_2991 = _zz_2992;
  assign _zz_2992 = ($signed(_zz_2993) >>> _zz_56);
  assign _zz_2993 = _zz_2994;
  assign _zz_2994 = ($signed(data_mid_26_real) + $signed(_zz_53));
  assign _zz_2995 = _zz_2996;
  assign _zz_2996 = ($signed(_zz_2997) >>> _zz_56);
  assign _zz_2997 = _zz_2998;
  assign _zz_2998 = ($signed(data_mid_26_imag) + $signed(_zz_54));
  assign _zz_2999 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_29_real));
  assign _zz_3000 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_29_imag));
  assign _zz_3001 = fixTo_28_dout;
  assign _zz_3002 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_29_imag));
  assign _zz_3003 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_29_real));
  assign _zz_3004 = fixTo_29_dout;
  assign _zz_3005 = _zz_3006;
  assign _zz_3006 = ($signed(_zz_3007) >>> _zz_59);
  assign _zz_3007 = _zz_3008;
  assign _zz_3008 = ($signed(data_mid_28_real) - $signed(_zz_57));
  assign _zz_3009 = _zz_3010;
  assign _zz_3010 = ($signed(_zz_3011) >>> _zz_59);
  assign _zz_3011 = _zz_3012;
  assign _zz_3012 = ($signed(data_mid_28_imag) - $signed(_zz_58));
  assign _zz_3013 = _zz_3014;
  assign _zz_3014 = ($signed(_zz_3015) >>> _zz_60);
  assign _zz_3015 = _zz_3016;
  assign _zz_3016 = ($signed(data_mid_28_real) + $signed(_zz_57));
  assign _zz_3017 = _zz_3018;
  assign _zz_3018 = ($signed(_zz_3019) >>> _zz_60);
  assign _zz_3019 = _zz_3020;
  assign _zz_3020 = ($signed(data_mid_28_imag) + $signed(_zz_58));
  assign _zz_3021 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_31_real));
  assign _zz_3022 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_31_imag));
  assign _zz_3023 = fixTo_30_dout;
  assign _zz_3024 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_31_imag));
  assign _zz_3025 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_31_real));
  assign _zz_3026 = fixTo_31_dout;
  assign _zz_3027 = _zz_3028;
  assign _zz_3028 = ($signed(_zz_3029) >>> _zz_63);
  assign _zz_3029 = _zz_3030;
  assign _zz_3030 = ($signed(data_mid_30_real) - $signed(_zz_61));
  assign _zz_3031 = _zz_3032;
  assign _zz_3032 = ($signed(_zz_3033) >>> _zz_63);
  assign _zz_3033 = _zz_3034;
  assign _zz_3034 = ($signed(data_mid_30_imag) - $signed(_zz_62));
  assign _zz_3035 = _zz_3036;
  assign _zz_3036 = ($signed(_zz_3037) >>> _zz_64);
  assign _zz_3037 = _zz_3038;
  assign _zz_3038 = ($signed(data_mid_30_real) + $signed(_zz_61));
  assign _zz_3039 = _zz_3040;
  assign _zz_3040 = ($signed(_zz_3041) >>> _zz_64);
  assign _zz_3041 = _zz_3042;
  assign _zz_3042 = ($signed(data_mid_30_imag) + $signed(_zz_62));
  assign _zz_3043 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_33_real));
  assign _zz_3044 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_33_imag));
  assign _zz_3045 = fixTo_32_dout;
  assign _zz_3046 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_33_imag));
  assign _zz_3047 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_33_real));
  assign _zz_3048 = fixTo_33_dout;
  assign _zz_3049 = _zz_3050;
  assign _zz_3050 = ($signed(_zz_3051) >>> _zz_67);
  assign _zz_3051 = _zz_3052;
  assign _zz_3052 = ($signed(data_mid_32_real) - $signed(_zz_65));
  assign _zz_3053 = _zz_3054;
  assign _zz_3054 = ($signed(_zz_3055) >>> _zz_67);
  assign _zz_3055 = _zz_3056;
  assign _zz_3056 = ($signed(data_mid_32_imag) - $signed(_zz_66));
  assign _zz_3057 = _zz_3058;
  assign _zz_3058 = ($signed(_zz_3059) >>> _zz_68);
  assign _zz_3059 = _zz_3060;
  assign _zz_3060 = ($signed(data_mid_32_real) + $signed(_zz_65));
  assign _zz_3061 = _zz_3062;
  assign _zz_3062 = ($signed(_zz_3063) >>> _zz_68);
  assign _zz_3063 = _zz_3064;
  assign _zz_3064 = ($signed(data_mid_32_imag) + $signed(_zz_66));
  assign _zz_3065 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_35_real));
  assign _zz_3066 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_35_imag));
  assign _zz_3067 = fixTo_34_dout;
  assign _zz_3068 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_35_imag));
  assign _zz_3069 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_35_real));
  assign _zz_3070 = fixTo_35_dout;
  assign _zz_3071 = _zz_3072;
  assign _zz_3072 = ($signed(_zz_3073) >>> _zz_71);
  assign _zz_3073 = _zz_3074;
  assign _zz_3074 = ($signed(data_mid_34_real) - $signed(_zz_69));
  assign _zz_3075 = _zz_3076;
  assign _zz_3076 = ($signed(_zz_3077) >>> _zz_71);
  assign _zz_3077 = _zz_3078;
  assign _zz_3078 = ($signed(data_mid_34_imag) - $signed(_zz_70));
  assign _zz_3079 = _zz_3080;
  assign _zz_3080 = ($signed(_zz_3081) >>> _zz_72);
  assign _zz_3081 = _zz_3082;
  assign _zz_3082 = ($signed(data_mid_34_real) + $signed(_zz_69));
  assign _zz_3083 = _zz_3084;
  assign _zz_3084 = ($signed(_zz_3085) >>> _zz_72);
  assign _zz_3085 = _zz_3086;
  assign _zz_3086 = ($signed(data_mid_34_imag) + $signed(_zz_70));
  assign _zz_3087 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_37_real));
  assign _zz_3088 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_37_imag));
  assign _zz_3089 = fixTo_36_dout;
  assign _zz_3090 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_37_imag));
  assign _zz_3091 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_37_real));
  assign _zz_3092 = fixTo_37_dout;
  assign _zz_3093 = _zz_3094;
  assign _zz_3094 = ($signed(_zz_3095) >>> _zz_75);
  assign _zz_3095 = _zz_3096;
  assign _zz_3096 = ($signed(data_mid_36_real) - $signed(_zz_73));
  assign _zz_3097 = _zz_3098;
  assign _zz_3098 = ($signed(_zz_3099) >>> _zz_75);
  assign _zz_3099 = _zz_3100;
  assign _zz_3100 = ($signed(data_mid_36_imag) - $signed(_zz_74));
  assign _zz_3101 = _zz_3102;
  assign _zz_3102 = ($signed(_zz_3103) >>> _zz_76);
  assign _zz_3103 = _zz_3104;
  assign _zz_3104 = ($signed(data_mid_36_real) + $signed(_zz_73));
  assign _zz_3105 = _zz_3106;
  assign _zz_3106 = ($signed(_zz_3107) >>> _zz_76);
  assign _zz_3107 = _zz_3108;
  assign _zz_3108 = ($signed(data_mid_36_imag) + $signed(_zz_74));
  assign _zz_3109 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_39_real));
  assign _zz_3110 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_39_imag));
  assign _zz_3111 = fixTo_38_dout;
  assign _zz_3112 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_39_imag));
  assign _zz_3113 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_39_real));
  assign _zz_3114 = fixTo_39_dout;
  assign _zz_3115 = _zz_3116;
  assign _zz_3116 = ($signed(_zz_3117) >>> _zz_79);
  assign _zz_3117 = _zz_3118;
  assign _zz_3118 = ($signed(data_mid_38_real) - $signed(_zz_77));
  assign _zz_3119 = _zz_3120;
  assign _zz_3120 = ($signed(_zz_3121) >>> _zz_79);
  assign _zz_3121 = _zz_3122;
  assign _zz_3122 = ($signed(data_mid_38_imag) - $signed(_zz_78));
  assign _zz_3123 = _zz_3124;
  assign _zz_3124 = ($signed(_zz_3125) >>> _zz_80);
  assign _zz_3125 = _zz_3126;
  assign _zz_3126 = ($signed(data_mid_38_real) + $signed(_zz_77));
  assign _zz_3127 = _zz_3128;
  assign _zz_3128 = ($signed(_zz_3129) >>> _zz_80);
  assign _zz_3129 = _zz_3130;
  assign _zz_3130 = ($signed(data_mid_38_imag) + $signed(_zz_78));
  assign _zz_3131 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_41_real));
  assign _zz_3132 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_41_imag));
  assign _zz_3133 = fixTo_40_dout;
  assign _zz_3134 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_41_imag));
  assign _zz_3135 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_41_real));
  assign _zz_3136 = fixTo_41_dout;
  assign _zz_3137 = _zz_3138;
  assign _zz_3138 = ($signed(_zz_3139) >>> _zz_83);
  assign _zz_3139 = _zz_3140;
  assign _zz_3140 = ($signed(data_mid_40_real) - $signed(_zz_81));
  assign _zz_3141 = _zz_3142;
  assign _zz_3142 = ($signed(_zz_3143) >>> _zz_83);
  assign _zz_3143 = _zz_3144;
  assign _zz_3144 = ($signed(data_mid_40_imag) - $signed(_zz_82));
  assign _zz_3145 = _zz_3146;
  assign _zz_3146 = ($signed(_zz_3147) >>> _zz_84);
  assign _zz_3147 = _zz_3148;
  assign _zz_3148 = ($signed(data_mid_40_real) + $signed(_zz_81));
  assign _zz_3149 = _zz_3150;
  assign _zz_3150 = ($signed(_zz_3151) >>> _zz_84);
  assign _zz_3151 = _zz_3152;
  assign _zz_3152 = ($signed(data_mid_40_imag) + $signed(_zz_82));
  assign _zz_3153 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_43_real));
  assign _zz_3154 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_43_imag));
  assign _zz_3155 = fixTo_42_dout;
  assign _zz_3156 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_43_imag));
  assign _zz_3157 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_43_real));
  assign _zz_3158 = fixTo_43_dout;
  assign _zz_3159 = _zz_3160;
  assign _zz_3160 = ($signed(_zz_3161) >>> _zz_87);
  assign _zz_3161 = _zz_3162;
  assign _zz_3162 = ($signed(data_mid_42_real) - $signed(_zz_85));
  assign _zz_3163 = _zz_3164;
  assign _zz_3164 = ($signed(_zz_3165) >>> _zz_87);
  assign _zz_3165 = _zz_3166;
  assign _zz_3166 = ($signed(data_mid_42_imag) - $signed(_zz_86));
  assign _zz_3167 = _zz_3168;
  assign _zz_3168 = ($signed(_zz_3169) >>> _zz_88);
  assign _zz_3169 = _zz_3170;
  assign _zz_3170 = ($signed(data_mid_42_real) + $signed(_zz_85));
  assign _zz_3171 = _zz_3172;
  assign _zz_3172 = ($signed(_zz_3173) >>> _zz_88);
  assign _zz_3173 = _zz_3174;
  assign _zz_3174 = ($signed(data_mid_42_imag) + $signed(_zz_86));
  assign _zz_3175 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_45_real));
  assign _zz_3176 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_45_imag));
  assign _zz_3177 = fixTo_44_dout;
  assign _zz_3178 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_45_imag));
  assign _zz_3179 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_45_real));
  assign _zz_3180 = fixTo_45_dout;
  assign _zz_3181 = _zz_3182;
  assign _zz_3182 = ($signed(_zz_3183) >>> _zz_91);
  assign _zz_3183 = _zz_3184;
  assign _zz_3184 = ($signed(data_mid_44_real) - $signed(_zz_89));
  assign _zz_3185 = _zz_3186;
  assign _zz_3186 = ($signed(_zz_3187) >>> _zz_91);
  assign _zz_3187 = _zz_3188;
  assign _zz_3188 = ($signed(data_mid_44_imag) - $signed(_zz_90));
  assign _zz_3189 = _zz_3190;
  assign _zz_3190 = ($signed(_zz_3191) >>> _zz_92);
  assign _zz_3191 = _zz_3192;
  assign _zz_3192 = ($signed(data_mid_44_real) + $signed(_zz_89));
  assign _zz_3193 = _zz_3194;
  assign _zz_3194 = ($signed(_zz_3195) >>> _zz_92);
  assign _zz_3195 = _zz_3196;
  assign _zz_3196 = ($signed(data_mid_44_imag) + $signed(_zz_90));
  assign _zz_3197 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_47_real));
  assign _zz_3198 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_47_imag));
  assign _zz_3199 = fixTo_46_dout;
  assign _zz_3200 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_47_imag));
  assign _zz_3201 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_47_real));
  assign _zz_3202 = fixTo_47_dout;
  assign _zz_3203 = _zz_3204;
  assign _zz_3204 = ($signed(_zz_3205) >>> _zz_95);
  assign _zz_3205 = _zz_3206;
  assign _zz_3206 = ($signed(data_mid_46_real) - $signed(_zz_93));
  assign _zz_3207 = _zz_3208;
  assign _zz_3208 = ($signed(_zz_3209) >>> _zz_95);
  assign _zz_3209 = _zz_3210;
  assign _zz_3210 = ($signed(data_mid_46_imag) - $signed(_zz_94));
  assign _zz_3211 = _zz_3212;
  assign _zz_3212 = ($signed(_zz_3213) >>> _zz_96);
  assign _zz_3213 = _zz_3214;
  assign _zz_3214 = ($signed(data_mid_46_real) + $signed(_zz_93));
  assign _zz_3215 = _zz_3216;
  assign _zz_3216 = ($signed(_zz_3217) >>> _zz_96);
  assign _zz_3217 = _zz_3218;
  assign _zz_3218 = ($signed(data_mid_46_imag) + $signed(_zz_94));
  assign _zz_3219 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_49_real));
  assign _zz_3220 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_49_imag));
  assign _zz_3221 = fixTo_48_dout;
  assign _zz_3222 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_49_imag));
  assign _zz_3223 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_49_real));
  assign _zz_3224 = fixTo_49_dout;
  assign _zz_3225 = _zz_3226;
  assign _zz_3226 = ($signed(_zz_3227) >>> _zz_99);
  assign _zz_3227 = _zz_3228;
  assign _zz_3228 = ($signed(data_mid_48_real) - $signed(_zz_97));
  assign _zz_3229 = _zz_3230;
  assign _zz_3230 = ($signed(_zz_3231) >>> _zz_99);
  assign _zz_3231 = _zz_3232;
  assign _zz_3232 = ($signed(data_mid_48_imag) - $signed(_zz_98));
  assign _zz_3233 = _zz_3234;
  assign _zz_3234 = ($signed(_zz_3235) >>> _zz_100);
  assign _zz_3235 = _zz_3236;
  assign _zz_3236 = ($signed(data_mid_48_real) + $signed(_zz_97));
  assign _zz_3237 = _zz_3238;
  assign _zz_3238 = ($signed(_zz_3239) >>> _zz_100);
  assign _zz_3239 = _zz_3240;
  assign _zz_3240 = ($signed(data_mid_48_imag) + $signed(_zz_98));
  assign _zz_3241 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_51_real));
  assign _zz_3242 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_51_imag));
  assign _zz_3243 = fixTo_50_dout;
  assign _zz_3244 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_51_imag));
  assign _zz_3245 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_51_real));
  assign _zz_3246 = fixTo_51_dout;
  assign _zz_3247 = _zz_3248;
  assign _zz_3248 = ($signed(_zz_3249) >>> _zz_103);
  assign _zz_3249 = _zz_3250;
  assign _zz_3250 = ($signed(data_mid_50_real) - $signed(_zz_101));
  assign _zz_3251 = _zz_3252;
  assign _zz_3252 = ($signed(_zz_3253) >>> _zz_103);
  assign _zz_3253 = _zz_3254;
  assign _zz_3254 = ($signed(data_mid_50_imag) - $signed(_zz_102));
  assign _zz_3255 = _zz_3256;
  assign _zz_3256 = ($signed(_zz_3257) >>> _zz_104);
  assign _zz_3257 = _zz_3258;
  assign _zz_3258 = ($signed(data_mid_50_real) + $signed(_zz_101));
  assign _zz_3259 = _zz_3260;
  assign _zz_3260 = ($signed(_zz_3261) >>> _zz_104);
  assign _zz_3261 = _zz_3262;
  assign _zz_3262 = ($signed(data_mid_50_imag) + $signed(_zz_102));
  assign _zz_3263 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_53_real));
  assign _zz_3264 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_53_imag));
  assign _zz_3265 = fixTo_52_dout;
  assign _zz_3266 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_53_imag));
  assign _zz_3267 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_53_real));
  assign _zz_3268 = fixTo_53_dout;
  assign _zz_3269 = _zz_3270;
  assign _zz_3270 = ($signed(_zz_3271) >>> _zz_107);
  assign _zz_3271 = _zz_3272;
  assign _zz_3272 = ($signed(data_mid_52_real) - $signed(_zz_105));
  assign _zz_3273 = _zz_3274;
  assign _zz_3274 = ($signed(_zz_3275) >>> _zz_107);
  assign _zz_3275 = _zz_3276;
  assign _zz_3276 = ($signed(data_mid_52_imag) - $signed(_zz_106));
  assign _zz_3277 = _zz_3278;
  assign _zz_3278 = ($signed(_zz_3279) >>> _zz_108);
  assign _zz_3279 = _zz_3280;
  assign _zz_3280 = ($signed(data_mid_52_real) + $signed(_zz_105));
  assign _zz_3281 = _zz_3282;
  assign _zz_3282 = ($signed(_zz_3283) >>> _zz_108);
  assign _zz_3283 = _zz_3284;
  assign _zz_3284 = ($signed(data_mid_52_imag) + $signed(_zz_106));
  assign _zz_3285 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_55_real));
  assign _zz_3286 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_55_imag));
  assign _zz_3287 = fixTo_54_dout;
  assign _zz_3288 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_55_imag));
  assign _zz_3289 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_55_real));
  assign _zz_3290 = fixTo_55_dout;
  assign _zz_3291 = _zz_3292;
  assign _zz_3292 = ($signed(_zz_3293) >>> _zz_111);
  assign _zz_3293 = _zz_3294;
  assign _zz_3294 = ($signed(data_mid_54_real) - $signed(_zz_109));
  assign _zz_3295 = _zz_3296;
  assign _zz_3296 = ($signed(_zz_3297) >>> _zz_111);
  assign _zz_3297 = _zz_3298;
  assign _zz_3298 = ($signed(data_mid_54_imag) - $signed(_zz_110));
  assign _zz_3299 = _zz_3300;
  assign _zz_3300 = ($signed(_zz_3301) >>> _zz_112);
  assign _zz_3301 = _zz_3302;
  assign _zz_3302 = ($signed(data_mid_54_real) + $signed(_zz_109));
  assign _zz_3303 = _zz_3304;
  assign _zz_3304 = ($signed(_zz_3305) >>> _zz_112);
  assign _zz_3305 = _zz_3306;
  assign _zz_3306 = ($signed(data_mid_54_imag) + $signed(_zz_110));
  assign _zz_3307 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_57_real));
  assign _zz_3308 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_57_imag));
  assign _zz_3309 = fixTo_56_dout;
  assign _zz_3310 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_57_imag));
  assign _zz_3311 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_57_real));
  assign _zz_3312 = fixTo_57_dout;
  assign _zz_3313 = _zz_3314;
  assign _zz_3314 = ($signed(_zz_3315) >>> _zz_115);
  assign _zz_3315 = _zz_3316;
  assign _zz_3316 = ($signed(data_mid_56_real) - $signed(_zz_113));
  assign _zz_3317 = _zz_3318;
  assign _zz_3318 = ($signed(_zz_3319) >>> _zz_115);
  assign _zz_3319 = _zz_3320;
  assign _zz_3320 = ($signed(data_mid_56_imag) - $signed(_zz_114));
  assign _zz_3321 = _zz_3322;
  assign _zz_3322 = ($signed(_zz_3323) >>> _zz_116);
  assign _zz_3323 = _zz_3324;
  assign _zz_3324 = ($signed(data_mid_56_real) + $signed(_zz_113));
  assign _zz_3325 = _zz_3326;
  assign _zz_3326 = ($signed(_zz_3327) >>> _zz_116);
  assign _zz_3327 = _zz_3328;
  assign _zz_3328 = ($signed(data_mid_56_imag) + $signed(_zz_114));
  assign _zz_3329 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_59_real));
  assign _zz_3330 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_59_imag));
  assign _zz_3331 = fixTo_58_dout;
  assign _zz_3332 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_59_imag));
  assign _zz_3333 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_59_real));
  assign _zz_3334 = fixTo_59_dout;
  assign _zz_3335 = _zz_3336;
  assign _zz_3336 = ($signed(_zz_3337) >>> _zz_119);
  assign _zz_3337 = _zz_3338;
  assign _zz_3338 = ($signed(data_mid_58_real) - $signed(_zz_117));
  assign _zz_3339 = _zz_3340;
  assign _zz_3340 = ($signed(_zz_3341) >>> _zz_119);
  assign _zz_3341 = _zz_3342;
  assign _zz_3342 = ($signed(data_mid_58_imag) - $signed(_zz_118));
  assign _zz_3343 = _zz_3344;
  assign _zz_3344 = ($signed(_zz_3345) >>> _zz_120);
  assign _zz_3345 = _zz_3346;
  assign _zz_3346 = ($signed(data_mid_58_real) + $signed(_zz_117));
  assign _zz_3347 = _zz_3348;
  assign _zz_3348 = ($signed(_zz_3349) >>> _zz_120);
  assign _zz_3349 = _zz_3350;
  assign _zz_3350 = ($signed(data_mid_58_imag) + $signed(_zz_118));
  assign _zz_3351 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_61_real));
  assign _zz_3352 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_61_imag));
  assign _zz_3353 = fixTo_60_dout;
  assign _zz_3354 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_61_imag));
  assign _zz_3355 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_61_real));
  assign _zz_3356 = fixTo_61_dout;
  assign _zz_3357 = _zz_3358;
  assign _zz_3358 = ($signed(_zz_3359) >>> _zz_123);
  assign _zz_3359 = _zz_3360;
  assign _zz_3360 = ($signed(data_mid_60_real) - $signed(_zz_121));
  assign _zz_3361 = _zz_3362;
  assign _zz_3362 = ($signed(_zz_3363) >>> _zz_123);
  assign _zz_3363 = _zz_3364;
  assign _zz_3364 = ($signed(data_mid_60_imag) - $signed(_zz_122));
  assign _zz_3365 = _zz_3366;
  assign _zz_3366 = ($signed(_zz_3367) >>> _zz_124);
  assign _zz_3367 = _zz_3368;
  assign _zz_3368 = ($signed(data_mid_60_real) + $signed(_zz_121));
  assign _zz_3369 = _zz_3370;
  assign _zz_3370 = ($signed(_zz_3371) >>> _zz_124);
  assign _zz_3371 = _zz_3372;
  assign _zz_3372 = ($signed(data_mid_60_imag) + $signed(_zz_122));
  assign _zz_3373 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_63_real));
  assign _zz_3374 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_63_imag));
  assign _zz_3375 = fixTo_62_dout;
  assign _zz_3376 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_63_imag));
  assign _zz_3377 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_63_real));
  assign _zz_3378 = fixTo_63_dout;
  assign _zz_3379 = _zz_3380;
  assign _zz_3380 = ($signed(_zz_3381) >>> _zz_127);
  assign _zz_3381 = _zz_3382;
  assign _zz_3382 = ($signed(data_mid_62_real) - $signed(_zz_125));
  assign _zz_3383 = _zz_3384;
  assign _zz_3384 = ($signed(_zz_3385) >>> _zz_127);
  assign _zz_3385 = _zz_3386;
  assign _zz_3386 = ($signed(data_mid_62_imag) - $signed(_zz_126));
  assign _zz_3387 = _zz_3388;
  assign _zz_3388 = ($signed(_zz_3389) >>> _zz_128);
  assign _zz_3389 = _zz_3390;
  assign _zz_3390 = ($signed(data_mid_62_real) + $signed(_zz_125));
  assign _zz_3391 = _zz_3392;
  assign _zz_3392 = ($signed(_zz_3393) >>> _zz_128);
  assign _zz_3393 = _zz_3394;
  assign _zz_3394 = ($signed(data_mid_62_imag) + $signed(_zz_126));
  assign _zz_3395 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_65_real));
  assign _zz_3396 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_65_imag));
  assign _zz_3397 = fixTo_64_dout;
  assign _zz_3398 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_65_imag));
  assign _zz_3399 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_65_real));
  assign _zz_3400 = fixTo_65_dout;
  assign _zz_3401 = _zz_3402;
  assign _zz_3402 = ($signed(_zz_3403) >>> _zz_131);
  assign _zz_3403 = _zz_3404;
  assign _zz_3404 = ($signed(data_mid_64_real) - $signed(_zz_129));
  assign _zz_3405 = _zz_3406;
  assign _zz_3406 = ($signed(_zz_3407) >>> _zz_131);
  assign _zz_3407 = _zz_3408;
  assign _zz_3408 = ($signed(data_mid_64_imag) - $signed(_zz_130));
  assign _zz_3409 = _zz_3410;
  assign _zz_3410 = ($signed(_zz_3411) >>> _zz_132);
  assign _zz_3411 = _zz_3412;
  assign _zz_3412 = ($signed(data_mid_64_real) + $signed(_zz_129));
  assign _zz_3413 = _zz_3414;
  assign _zz_3414 = ($signed(_zz_3415) >>> _zz_132);
  assign _zz_3415 = _zz_3416;
  assign _zz_3416 = ($signed(data_mid_64_imag) + $signed(_zz_130));
  assign _zz_3417 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_67_real));
  assign _zz_3418 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_67_imag));
  assign _zz_3419 = fixTo_66_dout;
  assign _zz_3420 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_67_imag));
  assign _zz_3421 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_67_real));
  assign _zz_3422 = fixTo_67_dout;
  assign _zz_3423 = _zz_3424;
  assign _zz_3424 = ($signed(_zz_3425) >>> _zz_135);
  assign _zz_3425 = _zz_3426;
  assign _zz_3426 = ($signed(data_mid_66_real) - $signed(_zz_133));
  assign _zz_3427 = _zz_3428;
  assign _zz_3428 = ($signed(_zz_3429) >>> _zz_135);
  assign _zz_3429 = _zz_3430;
  assign _zz_3430 = ($signed(data_mid_66_imag) - $signed(_zz_134));
  assign _zz_3431 = _zz_3432;
  assign _zz_3432 = ($signed(_zz_3433) >>> _zz_136);
  assign _zz_3433 = _zz_3434;
  assign _zz_3434 = ($signed(data_mid_66_real) + $signed(_zz_133));
  assign _zz_3435 = _zz_3436;
  assign _zz_3436 = ($signed(_zz_3437) >>> _zz_136);
  assign _zz_3437 = _zz_3438;
  assign _zz_3438 = ($signed(data_mid_66_imag) + $signed(_zz_134));
  assign _zz_3439 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_69_real));
  assign _zz_3440 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_69_imag));
  assign _zz_3441 = fixTo_68_dout;
  assign _zz_3442 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_69_imag));
  assign _zz_3443 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_69_real));
  assign _zz_3444 = fixTo_69_dout;
  assign _zz_3445 = _zz_3446;
  assign _zz_3446 = ($signed(_zz_3447) >>> _zz_139);
  assign _zz_3447 = _zz_3448;
  assign _zz_3448 = ($signed(data_mid_68_real) - $signed(_zz_137));
  assign _zz_3449 = _zz_3450;
  assign _zz_3450 = ($signed(_zz_3451) >>> _zz_139);
  assign _zz_3451 = _zz_3452;
  assign _zz_3452 = ($signed(data_mid_68_imag) - $signed(_zz_138));
  assign _zz_3453 = _zz_3454;
  assign _zz_3454 = ($signed(_zz_3455) >>> _zz_140);
  assign _zz_3455 = _zz_3456;
  assign _zz_3456 = ($signed(data_mid_68_real) + $signed(_zz_137));
  assign _zz_3457 = _zz_3458;
  assign _zz_3458 = ($signed(_zz_3459) >>> _zz_140);
  assign _zz_3459 = _zz_3460;
  assign _zz_3460 = ($signed(data_mid_68_imag) + $signed(_zz_138));
  assign _zz_3461 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_71_real));
  assign _zz_3462 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_71_imag));
  assign _zz_3463 = fixTo_70_dout;
  assign _zz_3464 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_71_imag));
  assign _zz_3465 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_71_real));
  assign _zz_3466 = fixTo_71_dout;
  assign _zz_3467 = _zz_3468;
  assign _zz_3468 = ($signed(_zz_3469) >>> _zz_143);
  assign _zz_3469 = _zz_3470;
  assign _zz_3470 = ($signed(data_mid_70_real) - $signed(_zz_141));
  assign _zz_3471 = _zz_3472;
  assign _zz_3472 = ($signed(_zz_3473) >>> _zz_143);
  assign _zz_3473 = _zz_3474;
  assign _zz_3474 = ($signed(data_mid_70_imag) - $signed(_zz_142));
  assign _zz_3475 = _zz_3476;
  assign _zz_3476 = ($signed(_zz_3477) >>> _zz_144);
  assign _zz_3477 = _zz_3478;
  assign _zz_3478 = ($signed(data_mid_70_real) + $signed(_zz_141));
  assign _zz_3479 = _zz_3480;
  assign _zz_3480 = ($signed(_zz_3481) >>> _zz_144);
  assign _zz_3481 = _zz_3482;
  assign _zz_3482 = ($signed(data_mid_70_imag) + $signed(_zz_142));
  assign _zz_3483 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_73_real));
  assign _zz_3484 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_73_imag));
  assign _zz_3485 = fixTo_72_dout;
  assign _zz_3486 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_73_imag));
  assign _zz_3487 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_73_real));
  assign _zz_3488 = fixTo_73_dout;
  assign _zz_3489 = _zz_3490;
  assign _zz_3490 = ($signed(_zz_3491) >>> _zz_147);
  assign _zz_3491 = _zz_3492;
  assign _zz_3492 = ($signed(data_mid_72_real) - $signed(_zz_145));
  assign _zz_3493 = _zz_3494;
  assign _zz_3494 = ($signed(_zz_3495) >>> _zz_147);
  assign _zz_3495 = _zz_3496;
  assign _zz_3496 = ($signed(data_mid_72_imag) - $signed(_zz_146));
  assign _zz_3497 = _zz_3498;
  assign _zz_3498 = ($signed(_zz_3499) >>> _zz_148);
  assign _zz_3499 = _zz_3500;
  assign _zz_3500 = ($signed(data_mid_72_real) + $signed(_zz_145));
  assign _zz_3501 = _zz_3502;
  assign _zz_3502 = ($signed(_zz_3503) >>> _zz_148);
  assign _zz_3503 = _zz_3504;
  assign _zz_3504 = ($signed(data_mid_72_imag) + $signed(_zz_146));
  assign _zz_3505 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_75_real));
  assign _zz_3506 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_75_imag));
  assign _zz_3507 = fixTo_74_dout;
  assign _zz_3508 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_75_imag));
  assign _zz_3509 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_75_real));
  assign _zz_3510 = fixTo_75_dout;
  assign _zz_3511 = _zz_3512;
  assign _zz_3512 = ($signed(_zz_3513) >>> _zz_151);
  assign _zz_3513 = _zz_3514;
  assign _zz_3514 = ($signed(data_mid_74_real) - $signed(_zz_149));
  assign _zz_3515 = _zz_3516;
  assign _zz_3516 = ($signed(_zz_3517) >>> _zz_151);
  assign _zz_3517 = _zz_3518;
  assign _zz_3518 = ($signed(data_mid_74_imag) - $signed(_zz_150));
  assign _zz_3519 = _zz_3520;
  assign _zz_3520 = ($signed(_zz_3521) >>> _zz_152);
  assign _zz_3521 = _zz_3522;
  assign _zz_3522 = ($signed(data_mid_74_real) + $signed(_zz_149));
  assign _zz_3523 = _zz_3524;
  assign _zz_3524 = ($signed(_zz_3525) >>> _zz_152);
  assign _zz_3525 = _zz_3526;
  assign _zz_3526 = ($signed(data_mid_74_imag) + $signed(_zz_150));
  assign _zz_3527 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_77_real));
  assign _zz_3528 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_77_imag));
  assign _zz_3529 = fixTo_76_dout;
  assign _zz_3530 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_77_imag));
  assign _zz_3531 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_77_real));
  assign _zz_3532 = fixTo_77_dout;
  assign _zz_3533 = _zz_3534;
  assign _zz_3534 = ($signed(_zz_3535) >>> _zz_155);
  assign _zz_3535 = _zz_3536;
  assign _zz_3536 = ($signed(data_mid_76_real) - $signed(_zz_153));
  assign _zz_3537 = _zz_3538;
  assign _zz_3538 = ($signed(_zz_3539) >>> _zz_155);
  assign _zz_3539 = _zz_3540;
  assign _zz_3540 = ($signed(data_mid_76_imag) - $signed(_zz_154));
  assign _zz_3541 = _zz_3542;
  assign _zz_3542 = ($signed(_zz_3543) >>> _zz_156);
  assign _zz_3543 = _zz_3544;
  assign _zz_3544 = ($signed(data_mid_76_real) + $signed(_zz_153));
  assign _zz_3545 = _zz_3546;
  assign _zz_3546 = ($signed(_zz_3547) >>> _zz_156);
  assign _zz_3547 = _zz_3548;
  assign _zz_3548 = ($signed(data_mid_76_imag) + $signed(_zz_154));
  assign _zz_3549 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_79_real));
  assign _zz_3550 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_79_imag));
  assign _zz_3551 = fixTo_78_dout;
  assign _zz_3552 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_79_imag));
  assign _zz_3553 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_79_real));
  assign _zz_3554 = fixTo_79_dout;
  assign _zz_3555 = _zz_3556;
  assign _zz_3556 = ($signed(_zz_3557) >>> _zz_159);
  assign _zz_3557 = _zz_3558;
  assign _zz_3558 = ($signed(data_mid_78_real) - $signed(_zz_157));
  assign _zz_3559 = _zz_3560;
  assign _zz_3560 = ($signed(_zz_3561) >>> _zz_159);
  assign _zz_3561 = _zz_3562;
  assign _zz_3562 = ($signed(data_mid_78_imag) - $signed(_zz_158));
  assign _zz_3563 = _zz_3564;
  assign _zz_3564 = ($signed(_zz_3565) >>> _zz_160);
  assign _zz_3565 = _zz_3566;
  assign _zz_3566 = ($signed(data_mid_78_real) + $signed(_zz_157));
  assign _zz_3567 = _zz_3568;
  assign _zz_3568 = ($signed(_zz_3569) >>> _zz_160);
  assign _zz_3569 = _zz_3570;
  assign _zz_3570 = ($signed(data_mid_78_imag) + $signed(_zz_158));
  assign _zz_3571 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_81_real));
  assign _zz_3572 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_81_imag));
  assign _zz_3573 = fixTo_80_dout;
  assign _zz_3574 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_81_imag));
  assign _zz_3575 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_81_real));
  assign _zz_3576 = fixTo_81_dout;
  assign _zz_3577 = _zz_3578;
  assign _zz_3578 = ($signed(_zz_3579) >>> _zz_163);
  assign _zz_3579 = _zz_3580;
  assign _zz_3580 = ($signed(data_mid_80_real) - $signed(_zz_161));
  assign _zz_3581 = _zz_3582;
  assign _zz_3582 = ($signed(_zz_3583) >>> _zz_163);
  assign _zz_3583 = _zz_3584;
  assign _zz_3584 = ($signed(data_mid_80_imag) - $signed(_zz_162));
  assign _zz_3585 = _zz_3586;
  assign _zz_3586 = ($signed(_zz_3587) >>> _zz_164);
  assign _zz_3587 = _zz_3588;
  assign _zz_3588 = ($signed(data_mid_80_real) + $signed(_zz_161));
  assign _zz_3589 = _zz_3590;
  assign _zz_3590 = ($signed(_zz_3591) >>> _zz_164);
  assign _zz_3591 = _zz_3592;
  assign _zz_3592 = ($signed(data_mid_80_imag) + $signed(_zz_162));
  assign _zz_3593 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_83_real));
  assign _zz_3594 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_83_imag));
  assign _zz_3595 = fixTo_82_dout;
  assign _zz_3596 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_83_imag));
  assign _zz_3597 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_83_real));
  assign _zz_3598 = fixTo_83_dout;
  assign _zz_3599 = _zz_3600;
  assign _zz_3600 = ($signed(_zz_3601) >>> _zz_167);
  assign _zz_3601 = _zz_3602;
  assign _zz_3602 = ($signed(data_mid_82_real) - $signed(_zz_165));
  assign _zz_3603 = _zz_3604;
  assign _zz_3604 = ($signed(_zz_3605) >>> _zz_167);
  assign _zz_3605 = _zz_3606;
  assign _zz_3606 = ($signed(data_mid_82_imag) - $signed(_zz_166));
  assign _zz_3607 = _zz_3608;
  assign _zz_3608 = ($signed(_zz_3609) >>> _zz_168);
  assign _zz_3609 = _zz_3610;
  assign _zz_3610 = ($signed(data_mid_82_real) + $signed(_zz_165));
  assign _zz_3611 = _zz_3612;
  assign _zz_3612 = ($signed(_zz_3613) >>> _zz_168);
  assign _zz_3613 = _zz_3614;
  assign _zz_3614 = ($signed(data_mid_82_imag) + $signed(_zz_166));
  assign _zz_3615 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_85_real));
  assign _zz_3616 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_85_imag));
  assign _zz_3617 = fixTo_84_dout;
  assign _zz_3618 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_85_imag));
  assign _zz_3619 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_85_real));
  assign _zz_3620 = fixTo_85_dout;
  assign _zz_3621 = _zz_3622;
  assign _zz_3622 = ($signed(_zz_3623) >>> _zz_171);
  assign _zz_3623 = _zz_3624;
  assign _zz_3624 = ($signed(data_mid_84_real) - $signed(_zz_169));
  assign _zz_3625 = _zz_3626;
  assign _zz_3626 = ($signed(_zz_3627) >>> _zz_171);
  assign _zz_3627 = _zz_3628;
  assign _zz_3628 = ($signed(data_mid_84_imag) - $signed(_zz_170));
  assign _zz_3629 = _zz_3630;
  assign _zz_3630 = ($signed(_zz_3631) >>> _zz_172);
  assign _zz_3631 = _zz_3632;
  assign _zz_3632 = ($signed(data_mid_84_real) + $signed(_zz_169));
  assign _zz_3633 = _zz_3634;
  assign _zz_3634 = ($signed(_zz_3635) >>> _zz_172);
  assign _zz_3635 = _zz_3636;
  assign _zz_3636 = ($signed(data_mid_84_imag) + $signed(_zz_170));
  assign _zz_3637 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_87_real));
  assign _zz_3638 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_87_imag));
  assign _zz_3639 = fixTo_86_dout;
  assign _zz_3640 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_87_imag));
  assign _zz_3641 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_87_real));
  assign _zz_3642 = fixTo_87_dout;
  assign _zz_3643 = _zz_3644;
  assign _zz_3644 = ($signed(_zz_3645) >>> _zz_175);
  assign _zz_3645 = _zz_3646;
  assign _zz_3646 = ($signed(data_mid_86_real) - $signed(_zz_173));
  assign _zz_3647 = _zz_3648;
  assign _zz_3648 = ($signed(_zz_3649) >>> _zz_175);
  assign _zz_3649 = _zz_3650;
  assign _zz_3650 = ($signed(data_mid_86_imag) - $signed(_zz_174));
  assign _zz_3651 = _zz_3652;
  assign _zz_3652 = ($signed(_zz_3653) >>> _zz_176);
  assign _zz_3653 = _zz_3654;
  assign _zz_3654 = ($signed(data_mid_86_real) + $signed(_zz_173));
  assign _zz_3655 = _zz_3656;
  assign _zz_3656 = ($signed(_zz_3657) >>> _zz_176);
  assign _zz_3657 = _zz_3658;
  assign _zz_3658 = ($signed(data_mid_86_imag) + $signed(_zz_174));
  assign _zz_3659 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_89_real));
  assign _zz_3660 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_89_imag));
  assign _zz_3661 = fixTo_88_dout;
  assign _zz_3662 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_89_imag));
  assign _zz_3663 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_89_real));
  assign _zz_3664 = fixTo_89_dout;
  assign _zz_3665 = _zz_3666;
  assign _zz_3666 = ($signed(_zz_3667) >>> _zz_179);
  assign _zz_3667 = _zz_3668;
  assign _zz_3668 = ($signed(data_mid_88_real) - $signed(_zz_177));
  assign _zz_3669 = _zz_3670;
  assign _zz_3670 = ($signed(_zz_3671) >>> _zz_179);
  assign _zz_3671 = _zz_3672;
  assign _zz_3672 = ($signed(data_mid_88_imag) - $signed(_zz_178));
  assign _zz_3673 = _zz_3674;
  assign _zz_3674 = ($signed(_zz_3675) >>> _zz_180);
  assign _zz_3675 = _zz_3676;
  assign _zz_3676 = ($signed(data_mid_88_real) + $signed(_zz_177));
  assign _zz_3677 = _zz_3678;
  assign _zz_3678 = ($signed(_zz_3679) >>> _zz_180);
  assign _zz_3679 = _zz_3680;
  assign _zz_3680 = ($signed(data_mid_88_imag) + $signed(_zz_178));
  assign _zz_3681 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_91_real));
  assign _zz_3682 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_91_imag));
  assign _zz_3683 = fixTo_90_dout;
  assign _zz_3684 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_91_imag));
  assign _zz_3685 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_91_real));
  assign _zz_3686 = fixTo_91_dout;
  assign _zz_3687 = _zz_3688;
  assign _zz_3688 = ($signed(_zz_3689) >>> _zz_183);
  assign _zz_3689 = _zz_3690;
  assign _zz_3690 = ($signed(data_mid_90_real) - $signed(_zz_181));
  assign _zz_3691 = _zz_3692;
  assign _zz_3692 = ($signed(_zz_3693) >>> _zz_183);
  assign _zz_3693 = _zz_3694;
  assign _zz_3694 = ($signed(data_mid_90_imag) - $signed(_zz_182));
  assign _zz_3695 = _zz_3696;
  assign _zz_3696 = ($signed(_zz_3697) >>> _zz_184);
  assign _zz_3697 = _zz_3698;
  assign _zz_3698 = ($signed(data_mid_90_real) + $signed(_zz_181));
  assign _zz_3699 = _zz_3700;
  assign _zz_3700 = ($signed(_zz_3701) >>> _zz_184);
  assign _zz_3701 = _zz_3702;
  assign _zz_3702 = ($signed(data_mid_90_imag) + $signed(_zz_182));
  assign _zz_3703 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_93_real));
  assign _zz_3704 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_93_imag));
  assign _zz_3705 = fixTo_92_dout;
  assign _zz_3706 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_93_imag));
  assign _zz_3707 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_93_real));
  assign _zz_3708 = fixTo_93_dout;
  assign _zz_3709 = _zz_3710;
  assign _zz_3710 = ($signed(_zz_3711) >>> _zz_187);
  assign _zz_3711 = _zz_3712;
  assign _zz_3712 = ($signed(data_mid_92_real) - $signed(_zz_185));
  assign _zz_3713 = _zz_3714;
  assign _zz_3714 = ($signed(_zz_3715) >>> _zz_187);
  assign _zz_3715 = _zz_3716;
  assign _zz_3716 = ($signed(data_mid_92_imag) - $signed(_zz_186));
  assign _zz_3717 = _zz_3718;
  assign _zz_3718 = ($signed(_zz_3719) >>> _zz_188);
  assign _zz_3719 = _zz_3720;
  assign _zz_3720 = ($signed(data_mid_92_real) + $signed(_zz_185));
  assign _zz_3721 = _zz_3722;
  assign _zz_3722 = ($signed(_zz_3723) >>> _zz_188);
  assign _zz_3723 = _zz_3724;
  assign _zz_3724 = ($signed(data_mid_92_imag) + $signed(_zz_186));
  assign _zz_3725 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_95_real));
  assign _zz_3726 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_95_imag));
  assign _zz_3727 = fixTo_94_dout;
  assign _zz_3728 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_95_imag));
  assign _zz_3729 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_95_real));
  assign _zz_3730 = fixTo_95_dout;
  assign _zz_3731 = _zz_3732;
  assign _zz_3732 = ($signed(_zz_3733) >>> _zz_191);
  assign _zz_3733 = _zz_3734;
  assign _zz_3734 = ($signed(data_mid_94_real) - $signed(_zz_189));
  assign _zz_3735 = _zz_3736;
  assign _zz_3736 = ($signed(_zz_3737) >>> _zz_191);
  assign _zz_3737 = _zz_3738;
  assign _zz_3738 = ($signed(data_mid_94_imag) - $signed(_zz_190));
  assign _zz_3739 = _zz_3740;
  assign _zz_3740 = ($signed(_zz_3741) >>> _zz_192);
  assign _zz_3741 = _zz_3742;
  assign _zz_3742 = ($signed(data_mid_94_real) + $signed(_zz_189));
  assign _zz_3743 = _zz_3744;
  assign _zz_3744 = ($signed(_zz_3745) >>> _zz_192);
  assign _zz_3745 = _zz_3746;
  assign _zz_3746 = ($signed(data_mid_94_imag) + $signed(_zz_190));
  assign _zz_3747 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_97_real));
  assign _zz_3748 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_97_imag));
  assign _zz_3749 = fixTo_96_dout;
  assign _zz_3750 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_97_imag));
  assign _zz_3751 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_97_real));
  assign _zz_3752 = fixTo_97_dout;
  assign _zz_3753 = _zz_3754;
  assign _zz_3754 = ($signed(_zz_3755) >>> _zz_195);
  assign _zz_3755 = _zz_3756;
  assign _zz_3756 = ($signed(data_mid_96_real) - $signed(_zz_193));
  assign _zz_3757 = _zz_3758;
  assign _zz_3758 = ($signed(_zz_3759) >>> _zz_195);
  assign _zz_3759 = _zz_3760;
  assign _zz_3760 = ($signed(data_mid_96_imag) - $signed(_zz_194));
  assign _zz_3761 = _zz_3762;
  assign _zz_3762 = ($signed(_zz_3763) >>> _zz_196);
  assign _zz_3763 = _zz_3764;
  assign _zz_3764 = ($signed(data_mid_96_real) + $signed(_zz_193));
  assign _zz_3765 = _zz_3766;
  assign _zz_3766 = ($signed(_zz_3767) >>> _zz_196);
  assign _zz_3767 = _zz_3768;
  assign _zz_3768 = ($signed(data_mid_96_imag) + $signed(_zz_194));
  assign _zz_3769 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_99_real));
  assign _zz_3770 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_99_imag));
  assign _zz_3771 = fixTo_98_dout;
  assign _zz_3772 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_99_imag));
  assign _zz_3773 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_99_real));
  assign _zz_3774 = fixTo_99_dout;
  assign _zz_3775 = _zz_3776;
  assign _zz_3776 = ($signed(_zz_3777) >>> _zz_199);
  assign _zz_3777 = _zz_3778;
  assign _zz_3778 = ($signed(data_mid_98_real) - $signed(_zz_197));
  assign _zz_3779 = _zz_3780;
  assign _zz_3780 = ($signed(_zz_3781) >>> _zz_199);
  assign _zz_3781 = _zz_3782;
  assign _zz_3782 = ($signed(data_mid_98_imag) - $signed(_zz_198));
  assign _zz_3783 = _zz_3784;
  assign _zz_3784 = ($signed(_zz_3785) >>> _zz_200);
  assign _zz_3785 = _zz_3786;
  assign _zz_3786 = ($signed(data_mid_98_real) + $signed(_zz_197));
  assign _zz_3787 = _zz_3788;
  assign _zz_3788 = ($signed(_zz_3789) >>> _zz_200);
  assign _zz_3789 = _zz_3790;
  assign _zz_3790 = ($signed(data_mid_98_imag) + $signed(_zz_198));
  assign _zz_3791 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_101_real));
  assign _zz_3792 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_101_imag));
  assign _zz_3793 = fixTo_100_dout;
  assign _zz_3794 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_101_imag));
  assign _zz_3795 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_101_real));
  assign _zz_3796 = fixTo_101_dout;
  assign _zz_3797 = _zz_3798;
  assign _zz_3798 = ($signed(_zz_3799) >>> _zz_203);
  assign _zz_3799 = _zz_3800;
  assign _zz_3800 = ($signed(data_mid_100_real) - $signed(_zz_201));
  assign _zz_3801 = _zz_3802;
  assign _zz_3802 = ($signed(_zz_3803) >>> _zz_203);
  assign _zz_3803 = _zz_3804;
  assign _zz_3804 = ($signed(data_mid_100_imag) - $signed(_zz_202));
  assign _zz_3805 = _zz_3806;
  assign _zz_3806 = ($signed(_zz_3807) >>> _zz_204);
  assign _zz_3807 = _zz_3808;
  assign _zz_3808 = ($signed(data_mid_100_real) + $signed(_zz_201));
  assign _zz_3809 = _zz_3810;
  assign _zz_3810 = ($signed(_zz_3811) >>> _zz_204);
  assign _zz_3811 = _zz_3812;
  assign _zz_3812 = ($signed(data_mid_100_imag) + $signed(_zz_202));
  assign _zz_3813 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_103_real));
  assign _zz_3814 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_103_imag));
  assign _zz_3815 = fixTo_102_dout;
  assign _zz_3816 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_103_imag));
  assign _zz_3817 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_103_real));
  assign _zz_3818 = fixTo_103_dout;
  assign _zz_3819 = _zz_3820;
  assign _zz_3820 = ($signed(_zz_3821) >>> _zz_207);
  assign _zz_3821 = _zz_3822;
  assign _zz_3822 = ($signed(data_mid_102_real) - $signed(_zz_205));
  assign _zz_3823 = _zz_3824;
  assign _zz_3824 = ($signed(_zz_3825) >>> _zz_207);
  assign _zz_3825 = _zz_3826;
  assign _zz_3826 = ($signed(data_mid_102_imag) - $signed(_zz_206));
  assign _zz_3827 = _zz_3828;
  assign _zz_3828 = ($signed(_zz_3829) >>> _zz_208);
  assign _zz_3829 = _zz_3830;
  assign _zz_3830 = ($signed(data_mid_102_real) + $signed(_zz_205));
  assign _zz_3831 = _zz_3832;
  assign _zz_3832 = ($signed(_zz_3833) >>> _zz_208);
  assign _zz_3833 = _zz_3834;
  assign _zz_3834 = ($signed(data_mid_102_imag) + $signed(_zz_206));
  assign _zz_3835 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_105_real));
  assign _zz_3836 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_105_imag));
  assign _zz_3837 = fixTo_104_dout;
  assign _zz_3838 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_105_imag));
  assign _zz_3839 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_105_real));
  assign _zz_3840 = fixTo_105_dout;
  assign _zz_3841 = _zz_3842;
  assign _zz_3842 = ($signed(_zz_3843) >>> _zz_211);
  assign _zz_3843 = _zz_3844;
  assign _zz_3844 = ($signed(data_mid_104_real) - $signed(_zz_209));
  assign _zz_3845 = _zz_3846;
  assign _zz_3846 = ($signed(_zz_3847) >>> _zz_211);
  assign _zz_3847 = _zz_3848;
  assign _zz_3848 = ($signed(data_mid_104_imag) - $signed(_zz_210));
  assign _zz_3849 = _zz_3850;
  assign _zz_3850 = ($signed(_zz_3851) >>> _zz_212);
  assign _zz_3851 = _zz_3852;
  assign _zz_3852 = ($signed(data_mid_104_real) + $signed(_zz_209));
  assign _zz_3853 = _zz_3854;
  assign _zz_3854 = ($signed(_zz_3855) >>> _zz_212);
  assign _zz_3855 = _zz_3856;
  assign _zz_3856 = ($signed(data_mid_104_imag) + $signed(_zz_210));
  assign _zz_3857 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_107_real));
  assign _zz_3858 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_107_imag));
  assign _zz_3859 = fixTo_106_dout;
  assign _zz_3860 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_107_imag));
  assign _zz_3861 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_107_real));
  assign _zz_3862 = fixTo_107_dout;
  assign _zz_3863 = _zz_3864;
  assign _zz_3864 = ($signed(_zz_3865) >>> _zz_215);
  assign _zz_3865 = _zz_3866;
  assign _zz_3866 = ($signed(data_mid_106_real) - $signed(_zz_213));
  assign _zz_3867 = _zz_3868;
  assign _zz_3868 = ($signed(_zz_3869) >>> _zz_215);
  assign _zz_3869 = _zz_3870;
  assign _zz_3870 = ($signed(data_mid_106_imag) - $signed(_zz_214));
  assign _zz_3871 = _zz_3872;
  assign _zz_3872 = ($signed(_zz_3873) >>> _zz_216);
  assign _zz_3873 = _zz_3874;
  assign _zz_3874 = ($signed(data_mid_106_real) + $signed(_zz_213));
  assign _zz_3875 = _zz_3876;
  assign _zz_3876 = ($signed(_zz_3877) >>> _zz_216);
  assign _zz_3877 = _zz_3878;
  assign _zz_3878 = ($signed(data_mid_106_imag) + $signed(_zz_214));
  assign _zz_3879 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_109_real));
  assign _zz_3880 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_109_imag));
  assign _zz_3881 = fixTo_108_dout;
  assign _zz_3882 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_109_imag));
  assign _zz_3883 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_109_real));
  assign _zz_3884 = fixTo_109_dout;
  assign _zz_3885 = _zz_3886;
  assign _zz_3886 = ($signed(_zz_3887) >>> _zz_219);
  assign _zz_3887 = _zz_3888;
  assign _zz_3888 = ($signed(data_mid_108_real) - $signed(_zz_217));
  assign _zz_3889 = _zz_3890;
  assign _zz_3890 = ($signed(_zz_3891) >>> _zz_219);
  assign _zz_3891 = _zz_3892;
  assign _zz_3892 = ($signed(data_mid_108_imag) - $signed(_zz_218));
  assign _zz_3893 = _zz_3894;
  assign _zz_3894 = ($signed(_zz_3895) >>> _zz_220);
  assign _zz_3895 = _zz_3896;
  assign _zz_3896 = ($signed(data_mid_108_real) + $signed(_zz_217));
  assign _zz_3897 = _zz_3898;
  assign _zz_3898 = ($signed(_zz_3899) >>> _zz_220);
  assign _zz_3899 = _zz_3900;
  assign _zz_3900 = ($signed(data_mid_108_imag) + $signed(_zz_218));
  assign _zz_3901 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_111_real));
  assign _zz_3902 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_111_imag));
  assign _zz_3903 = fixTo_110_dout;
  assign _zz_3904 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_111_imag));
  assign _zz_3905 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_111_real));
  assign _zz_3906 = fixTo_111_dout;
  assign _zz_3907 = _zz_3908;
  assign _zz_3908 = ($signed(_zz_3909) >>> _zz_223);
  assign _zz_3909 = _zz_3910;
  assign _zz_3910 = ($signed(data_mid_110_real) - $signed(_zz_221));
  assign _zz_3911 = _zz_3912;
  assign _zz_3912 = ($signed(_zz_3913) >>> _zz_223);
  assign _zz_3913 = _zz_3914;
  assign _zz_3914 = ($signed(data_mid_110_imag) - $signed(_zz_222));
  assign _zz_3915 = _zz_3916;
  assign _zz_3916 = ($signed(_zz_3917) >>> _zz_224);
  assign _zz_3917 = _zz_3918;
  assign _zz_3918 = ($signed(data_mid_110_real) + $signed(_zz_221));
  assign _zz_3919 = _zz_3920;
  assign _zz_3920 = ($signed(_zz_3921) >>> _zz_224);
  assign _zz_3921 = _zz_3922;
  assign _zz_3922 = ($signed(data_mid_110_imag) + $signed(_zz_222));
  assign _zz_3923 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_113_real));
  assign _zz_3924 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_113_imag));
  assign _zz_3925 = fixTo_112_dout;
  assign _zz_3926 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_113_imag));
  assign _zz_3927 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_113_real));
  assign _zz_3928 = fixTo_113_dout;
  assign _zz_3929 = _zz_3930;
  assign _zz_3930 = ($signed(_zz_3931) >>> _zz_227);
  assign _zz_3931 = _zz_3932;
  assign _zz_3932 = ($signed(data_mid_112_real) - $signed(_zz_225));
  assign _zz_3933 = _zz_3934;
  assign _zz_3934 = ($signed(_zz_3935) >>> _zz_227);
  assign _zz_3935 = _zz_3936;
  assign _zz_3936 = ($signed(data_mid_112_imag) - $signed(_zz_226));
  assign _zz_3937 = _zz_3938;
  assign _zz_3938 = ($signed(_zz_3939) >>> _zz_228);
  assign _zz_3939 = _zz_3940;
  assign _zz_3940 = ($signed(data_mid_112_real) + $signed(_zz_225));
  assign _zz_3941 = _zz_3942;
  assign _zz_3942 = ($signed(_zz_3943) >>> _zz_228);
  assign _zz_3943 = _zz_3944;
  assign _zz_3944 = ($signed(data_mid_112_imag) + $signed(_zz_226));
  assign _zz_3945 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_115_real));
  assign _zz_3946 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_115_imag));
  assign _zz_3947 = fixTo_114_dout;
  assign _zz_3948 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_115_imag));
  assign _zz_3949 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_115_real));
  assign _zz_3950 = fixTo_115_dout;
  assign _zz_3951 = _zz_3952;
  assign _zz_3952 = ($signed(_zz_3953) >>> _zz_231);
  assign _zz_3953 = _zz_3954;
  assign _zz_3954 = ($signed(data_mid_114_real) - $signed(_zz_229));
  assign _zz_3955 = _zz_3956;
  assign _zz_3956 = ($signed(_zz_3957) >>> _zz_231);
  assign _zz_3957 = _zz_3958;
  assign _zz_3958 = ($signed(data_mid_114_imag) - $signed(_zz_230));
  assign _zz_3959 = _zz_3960;
  assign _zz_3960 = ($signed(_zz_3961) >>> _zz_232);
  assign _zz_3961 = _zz_3962;
  assign _zz_3962 = ($signed(data_mid_114_real) + $signed(_zz_229));
  assign _zz_3963 = _zz_3964;
  assign _zz_3964 = ($signed(_zz_3965) >>> _zz_232);
  assign _zz_3965 = _zz_3966;
  assign _zz_3966 = ($signed(data_mid_114_imag) + $signed(_zz_230));
  assign _zz_3967 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_117_real));
  assign _zz_3968 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_117_imag));
  assign _zz_3969 = fixTo_116_dout;
  assign _zz_3970 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_117_imag));
  assign _zz_3971 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_117_real));
  assign _zz_3972 = fixTo_117_dout;
  assign _zz_3973 = _zz_3974;
  assign _zz_3974 = ($signed(_zz_3975) >>> _zz_235);
  assign _zz_3975 = _zz_3976;
  assign _zz_3976 = ($signed(data_mid_116_real) - $signed(_zz_233));
  assign _zz_3977 = _zz_3978;
  assign _zz_3978 = ($signed(_zz_3979) >>> _zz_235);
  assign _zz_3979 = _zz_3980;
  assign _zz_3980 = ($signed(data_mid_116_imag) - $signed(_zz_234));
  assign _zz_3981 = _zz_3982;
  assign _zz_3982 = ($signed(_zz_3983) >>> _zz_236);
  assign _zz_3983 = _zz_3984;
  assign _zz_3984 = ($signed(data_mid_116_real) + $signed(_zz_233));
  assign _zz_3985 = _zz_3986;
  assign _zz_3986 = ($signed(_zz_3987) >>> _zz_236);
  assign _zz_3987 = _zz_3988;
  assign _zz_3988 = ($signed(data_mid_116_imag) + $signed(_zz_234));
  assign _zz_3989 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_119_real));
  assign _zz_3990 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_119_imag));
  assign _zz_3991 = fixTo_118_dout;
  assign _zz_3992 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_119_imag));
  assign _zz_3993 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_119_real));
  assign _zz_3994 = fixTo_119_dout;
  assign _zz_3995 = _zz_3996;
  assign _zz_3996 = ($signed(_zz_3997) >>> _zz_239);
  assign _zz_3997 = _zz_3998;
  assign _zz_3998 = ($signed(data_mid_118_real) - $signed(_zz_237));
  assign _zz_3999 = _zz_4000;
  assign _zz_4000 = ($signed(_zz_4001) >>> _zz_239);
  assign _zz_4001 = _zz_4002;
  assign _zz_4002 = ($signed(data_mid_118_imag) - $signed(_zz_238));
  assign _zz_4003 = _zz_4004;
  assign _zz_4004 = ($signed(_zz_4005) >>> _zz_240);
  assign _zz_4005 = _zz_4006;
  assign _zz_4006 = ($signed(data_mid_118_real) + $signed(_zz_237));
  assign _zz_4007 = _zz_4008;
  assign _zz_4008 = ($signed(_zz_4009) >>> _zz_240);
  assign _zz_4009 = _zz_4010;
  assign _zz_4010 = ($signed(data_mid_118_imag) + $signed(_zz_238));
  assign _zz_4011 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_121_real));
  assign _zz_4012 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_121_imag));
  assign _zz_4013 = fixTo_120_dout;
  assign _zz_4014 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_121_imag));
  assign _zz_4015 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_121_real));
  assign _zz_4016 = fixTo_121_dout;
  assign _zz_4017 = _zz_4018;
  assign _zz_4018 = ($signed(_zz_4019) >>> _zz_243);
  assign _zz_4019 = _zz_4020;
  assign _zz_4020 = ($signed(data_mid_120_real) - $signed(_zz_241));
  assign _zz_4021 = _zz_4022;
  assign _zz_4022 = ($signed(_zz_4023) >>> _zz_243);
  assign _zz_4023 = _zz_4024;
  assign _zz_4024 = ($signed(data_mid_120_imag) - $signed(_zz_242));
  assign _zz_4025 = _zz_4026;
  assign _zz_4026 = ($signed(_zz_4027) >>> _zz_244);
  assign _zz_4027 = _zz_4028;
  assign _zz_4028 = ($signed(data_mid_120_real) + $signed(_zz_241));
  assign _zz_4029 = _zz_4030;
  assign _zz_4030 = ($signed(_zz_4031) >>> _zz_244);
  assign _zz_4031 = _zz_4032;
  assign _zz_4032 = ($signed(data_mid_120_imag) + $signed(_zz_242));
  assign _zz_4033 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_123_real));
  assign _zz_4034 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_123_imag));
  assign _zz_4035 = fixTo_122_dout;
  assign _zz_4036 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_123_imag));
  assign _zz_4037 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_123_real));
  assign _zz_4038 = fixTo_123_dout;
  assign _zz_4039 = _zz_4040;
  assign _zz_4040 = ($signed(_zz_4041) >>> _zz_247);
  assign _zz_4041 = _zz_4042;
  assign _zz_4042 = ($signed(data_mid_122_real) - $signed(_zz_245));
  assign _zz_4043 = _zz_4044;
  assign _zz_4044 = ($signed(_zz_4045) >>> _zz_247);
  assign _zz_4045 = _zz_4046;
  assign _zz_4046 = ($signed(data_mid_122_imag) - $signed(_zz_246));
  assign _zz_4047 = _zz_4048;
  assign _zz_4048 = ($signed(_zz_4049) >>> _zz_248);
  assign _zz_4049 = _zz_4050;
  assign _zz_4050 = ($signed(data_mid_122_real) + $signed(_zz_245));
  assign _zz_4051 = _zz_4052;
  assign _zz_4052 = ($signed(_zz_4053) >>> _zz_248);
  assign _zz_4053 = _zz_4054;
  assign _zz_4054 = ($signed(data_mid_122_imag) + $signed(_zz_246));
  assign _zz_4055 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_125_real));
  assign _zz_4056 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_125_imag));
  assign _zz_4057 = fixTo_124_dout;
  assign _zz_4058 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_125_imag));
  assign _zz_4059 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_125_real));
  assign _zz_4060 = fixTo_125_dout;
  assign _zz_4061 = _zz_4062;
  assign _zz_4062 = ($signed(_zz_4063) >>> _zz_251);
  assign _zz_4063 = _zz_4064;
  assign _zz_4064 = ($signed(data_mid_124_real) - $signed(_zz_249));
  assign _zz_4065 = _zz_4066;
  assign _zz_4066 = ($signed(_zz_4067) >>> _zz_251);
  assign _zz_4067 = _zz_4068;
  assign _zz_4068 = ($signed(data_mid_124_imag) - $signed(_zz_250));
  assign _zz_4069 = _zz_4070;
  assign _zz_4070 = ($signed(_zz_4071) >>> _zz_252);
  assign _zz_4071 = _zz_4072;
  assign _zz_4072 = ($signed(data_mid_124_real) + $signed(_zz_249));
  assign _zz_4073 = _zz_4074;
  assign _zz_4074 = ($signed(_zz_4075) >>> _zz_252);
  assign _zz_4075 = _zz_4076;
  assign _zz_4076 = ($signed(data_mid_124_imag) + $signed(_zz_250));
  assign _zz_4077 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_127_real));
  assign _zz_4078 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_127_imag));
  assign _zz_4079 = fixTo_126_dout;
  assign _zz_4080 = ($signed(twiddle_factor_table_0_real) * $signed(data_mid_127_imag));
  assign _zz_4081 = ($signed(twiddle_factor_table_0_imag) * $signed(data_mid_127_real));
  assign _zz_4082 = fixTo_127_dout;
  assign _zz_4083 = _zz_4084;
  assign _zz_4084 = ($signed(_zz_4085) >>> _zz_255);
  assign _zz_4085 = _zz_4086;
  assign _zz_4086 = ($signed(data_mid_126_real) - $signed(_zz_253));
  assign _zz_4087 = _zz_4088;
  assign _zz_4088 = ($signed(_zz_4089) >>> _zz_255);
  assign _zz_4089 = _zz_4090;
  assign _zz_4090 = ($signed(data_mid_126_imag) - $signed(_zz_254));
  assign _zz_4091 = _zz_4092;
  assign _zz_4092 = ($signed(_zz_4093) >>> _zz_256);
  assign _zz_4093 = _zz_4094;
  assign _zz_4094 = ($signed(data_mid_126_real) + $signed(_zz_253));
  assign _zz_4095 = _zz_4096;
  assign _zz_4096 = ($signed(_zz_4097) >>> _zz_256);
  assign _zz_4097 = _zz_4098;
  assign _zz_4098 = ($signed(data_mid_126_imag) + $signed(_zz_254));
  assign _zz_4099 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_2_real));
  assign _zz_4100 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_2_imag));
  assign _zz_4101 = fixTo_128_dout;
  assign _zz_4102 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_2_imag));
  assign _zz_4103 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_2_real));
  assign _zz_4104 = fixTo_129_dout;
  assign _zz_4105 = _zz_4106;
  assign _zz_4106 = ($signed(_zz_4107) >>> _zz_259);
  assign _zz_4107 = _zz_4108;
  assign _zz_4108 = ($signed(data_mid_0_real) - $signed(_zz_257));
  assign _zz_4109 = _zz_4110;
  assign _zz_4110 = ($signed(_zz_4111) >>> _zz_259);
  assign _zz_4111 = _zz_4112;
  assign _zz_4112 = ($signed(data_mid_0_imag) - $signed(_zz_258));
  assign _zz_4113 = _zz_4114;
  assign _zz_4114 = ($signed(_zz_4115) >>> _zz_260);
  assign _zz_4115 = _zz_4116;
  assign _zz_4116 = ($signed(data_mid_0_real) + $signed(_zz_257));
  assign _zz_4117 = _zz_4118;
  assign _zz_4118 = ($signed(_zz_4119) >>> _zz_260);
  assign _zz_4119 = _zz_4120;
  assign _zz_4120 = ($signed(data_mid_0_imag) + $signed(_zz_258));
  assign _zz_4121 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_3_real));
  assign _zz_4122 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_3_imag));
  assign _zz_4123 = fixTo_130_dout;
  assign _zz_4124 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_3_imag));
  assign _zz_4125 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_3_real));
  assign _zz_4126 = fixTo_131_dout;
  assign _zz_4127 = _zz_4128;
  assign _zz_4128 = ($signed(_zz_4129) >>> _zz_263);
  assign _zz_4129 = _zz_4130;
  assign _zz_4130 = ($signed(data_mid_1_real) - $signed(_zz_261));
  assign _zz_4131 = _zz_4132;
  assign _zz_4132 = ($signed(_zz_4133) >>> _zz_263);
  assign _zz_4133 = _zz_4134;
  assign _zz_4134 = ($signed(data_mid_1_imag) - $signed(_zz_262));
  assign _zz_4135 = _zz_4136;
  assign _zz_4136 = ($signed(_zz_4137) >>> _zz_264);
  assign _zz_4137 = _zz_4138;
  assign _zz_4138 = ($signed(data_mid_1_real) + $signed(_zz_261));
  assign _zz_4139 = _zz_4140;
  assign _zz_4140 = ($signed(_zz_4141) >>> _zz_264);
  assign _zz_4141 = _zz_4142;
  assign _zz_4142 = ($signed(data_mid_1_imag) + $signed(_zz_262));
  assign _zz_4143 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_6_real));
  assign _zz_4144 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_6_imag));
  assign _zz_4145 = fixTo_132_dout;
  assign _zz_4146 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_6_imag));
  assign _zz_4147 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_6_real));
  assign _zz_4148 = fixTo_133_dout;
  assign _zz_4149 = _zz_4150;
  assign _zz_4150 = ($signed(_zz_4151) >>> _zz_267);
  assign _zz_4151 = _zz_4152;
  assign _zz_4152 = ($signed(data_mid_4_real) - $signed(_zz_265));
  assign _zz_4153 = _zz_4154;
  assign _zz_4154 = ($signed(_zz_4155) >>> _zz_267);
  assign _zz_4155 = _zz_4156;
  assign _zz_4156 = ($signed(data_mid_4_imag) - $signed(_zz_266));
  assign _zz_4157 = _zz_4158;
  assign _zz_4158 = ($signed(_zz_4159) >>> _zz_268);
  assign _zz_4159 = _zz_4160;
  assign _zz_4160 = ($signed(data_mid_4_real) + $signed(_zz_265));
  assign _zz_4161 = _zz_4162;
  assign _zz_4162 = ($signed(_zz_4163) >>> _zz_268);
  assign _zz_4163 = _zz_4164;
  assign _zz_4164 = ($signed(data_mid_4_imag) + $signed(_zz_266));
  assign _zz_4165 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_7_real));
  assign _zz_4166 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_7_imag));
  assign _zz_4167 = fixTo_134_dout;
  assign _zz_4168 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_7_imag));
  assign _zz_4169 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_7_real));
  assign _zz_4170 = fixTo_135_dout;
  assign _zz_4171 = _zz_4172;
  assign _zz_4172 = ($signed(_zz_4173) >>> _zz_271);
  assign _zz_4173 = _zz_4174;
  assign _zz_4174 = ($signed(data_mid_5_real) - $signed(_zz_269));
  assign _zz_4175 = _zz_4176;
  assign _zz_4176 = ($signed(_zz_4177) >>> _zz_271);
  assign _zz_4177 = _zz_4178;
  assign _zz_4178 = ($signed(data_mid_5_imag) - $signed(_zz_270));
  assign _zz_4179 = _zz_4180;
  assign _zz_4180 = ($signed(_zz_4181) >>> _zz_272);
  assign _zz_4181 = _zz_4182;
  assign _zz_4182 = ($signed(data_mid_5_real) + $signed(_zz_269));
  assign _zz_4183 = _zz_4184;
  assign _zz_4184 = ($signed(_zz_4185) >>> _zz_272);
  assign _zz_4185 = _zz_4186;
  assign _zz_4186 = ($signed(data_mid_5_imag) + $signed(_zz_270));
  assign _zz_4187 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_10_real));
  assign _zz_4188 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_10_imag));
  assign _zz_4189 = fixTo_136_dout;
  assign _zz_4190 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_10_imag));
  assign _zz_4191 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_10_real));
  assign _zz_4192 = fixTo_137_dout;
  assign _zz_4193 = _zz_4194;
  assign _zz_4194 = ($signed(_zz_4195) >>> _zz_275);
  assign _zz_4195 = _zz_4196;
  assign _zz_4196 = ($signed(data_mid_8_real) - $signed(_zz_273));
  assign _zz_4197 = _zz_4198;
  assign _zz_4198 = ($signed(_zz_4199) >>> _zz_275);
  assign _zz_4199 = _zz_4200;
  assign _zz_4200 = ($signed(data_mid_8_imag) - $signed(_zz_274));
  assign _zz_4201 = _zz_4202;
  assign _zz_4202 = ($signed(_zz_4203) >>> _zz_276);
  assign _zz_4203 = _zz_4204;
  assign _zz_4204 = ($signed(data_mid_8_real) + $signed(_zz_273));
  assign _zz_4205 = _zz_4206;
  assign _zz_4206 = ($signed(_zz_4207) >>> _zz_276);
  assign _zz_4207 = _zz_4208;
  assign _zz_4208 = ($signed(data_mid_8_imag) + $signed(_zz_274));
  assign _zz_4209 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_11_real));
  assign _zz_4210 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_11_imag));
  assign _zz_4211 = fixTo_138_dout;
  assign _zz_4212 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_11_imag));
  assign _zz_4213 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_11_real));
  assign _zz_4214 = fixTo_139_dout;
  assign _zz_4215 = _zz_4216;
  assign _zz_4216 = ($signed(_zz_4217) >>> _zz_279);
  assign _zz_4217 = _zz_4218;
  assign _zz_4218 = ($signed(data_mid_9_real) - $signed(_zz_277));
  assign _zz_4219 = _zz_4220;
  assign _zz_4220 = ($signed(_zz_4221) >>> _zz_279);
  assign _zz_4221 = _zz_4222;
  assign _zz_4222 = ($signed(data_mid_9_imag) - $signed(_zz_278));
  assign _zz_4223 = _zz_4224;
  assign _zz_4224 = ($signed(_zz_4225) >>> _zz_280);
  assign _zz_4225 = _zz_4226;
  assign _zz_4226 = ($signed(data_mid_9_real) + $signed(_zz_277));
  assign _zz_4227 = _zz_4228;
  assign _zz_4228 = ($signed(_zz_4229) >>> _zz_280);
  assign _zz_4229 = _zz_4230;
  assign _zz_4230 = ($signed(data_mid_9_imag) + $signed(_zz_278));
  assign _zz_4231 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_14_real));
  assign _zz_4232 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_14_imag));
  assign _zz_4233 = fixTo_140_dout;
  assign _zz_4234 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_14_imag));
  assign _zz_4235 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_14_real));
  assign _zz_4236 = fixTo_141_dout;
  assign _zz_4237 = _zz_4238;
  assign _zz_4238 = ($signed(_zz_4239) >>> _zz_283);
  assign _zz_4239 = _zz_4240;
  assign _zz_4240 = ($signed(data_mid_12_real) - $signed(_zz_281));
  assign _zz_4241 = _zz_4242;
  assign _zz_4242 = ($signed(_zz_4243) >>> _zz_283);
  assign _zz_4243 = _zz_4244;
  assign _zz_4244 = ($signed(data_mid_12_imag) - $signed(_zz_282));
  assign _zz_4245 = _zz_4246;
  assign _zz_4246 = ($signed(_zz_4247) >>> _zz_284);
  assign _zz_4247 = _zz_4248;
  assign _zz_4248 = ($signed(data_mid_12_real) + $signed(_zz_281));
  assign _zz_4249 = _zz_4250;
  assign _zz_4250 = ($signed(_zz_4251) >>> _zz_284);
  assign _zz_4251 = _zz_4252;
  assign _zz_4252 = ($signed(data_mid_12_imag) + $signed(_zz_282));
  assign _zz_4253 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_15_real));
  assign _zz_4254 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_15_imag));
  assign _zz_4255 = fixTo_142_dout;
  assign _zz_4256 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_15_imag));
  assign _zz_4257 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_15_real));
  assign _zz_4258 = fixTo_143_dout;
  assign _zz_4259 = _zz_4260;
  assign _zz_4260 = ($signed(_zz_4261) >>> _zz_287);
  assign _zz_4261 = _zz_4262;
  assign _zz_4262 = ($signed(data_mid_13_real) - $signed(_zz_285));
  assign _zz_4263 = _zz_4264;
  assign _zz_4264 = ($signed(_zz_4265) >>> _zz_287);
  assign _zz_4265 = _zz_4266;
  assign _zz_4266 = ($signed(data_mid_13_imag) - $signed(_zz_286));
  assign _zz_4267 = _zz_4268;
  assign _zz_4268 = ($signed(_zz_4269) >>> _zz_288);
  assign _zz_4269 = _zz_4270;
  assign _zz_4270 = ($signed(data_mid_13_real) + $signed(_zz_285));
  assign _zz_4271 = _zz_4272;
  assign _zz_4272 = ($signed(_zz_4273) >>> _zz_288);
  assign _zz_4273 = _zz_4274;
  assign _zz_4274 = ($signed(data_mid_13_imag) + $signed(_zz_286));
  assign _zz_4275 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_18_real));
  assign _zz_4276 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_18_imag));
  assign _zz_4277 = fixTo_144_dout;
  assign _zz_4278 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_18_imag));
  assign _zz_4279 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_18_real));
  assign _zz_4280 = fixTo_145_dout;
  assign _zz_4281 = _zz_4282;
  assign _zz_4282 = ($signed(_zz_4283) >>> _zz_291);
  assign _zz_4283 = _zz_4284;
  assign _zz_4284 = ($signed(data_mid_16_real) - $signed(_zz_289));
  assign _zz_4285 = _zz_4286;
  assign _zz_4286 = ($signed(_zz_4287) >>> _zz_291);
  assign _zz_4287 = _zz_4288;
  assign _zz_4288 = ($signed(data_mid_16_imag) - $signed(_zz_290));
  assign _zz_4289 = _zz_4290;
  assign _zz_4290 = ($signed(_zz_4291) >>> _zz_292);
  assign _zz_4291 = _zz_4292;
  assign _zz_4292 = ($signed(data_mid_16_real) + $signed(_zz_289));
  assign _zz_4293 = _zz_4294;
  assign _zz_4294 = ($signed(_zz_4295) >>> _zz_292);
  assign _zz_4295 = _zz_4296;
  assign _zz_4296 = ($signed(data_mid_16_imag) + $signed(_zz_290));
  assign _zz_4297 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_19_real));
  assign _zz_4298 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_19_imag));
  assign _zz_4299 = fixTo_146_dout;
  assign _zz_4300 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_19_imag));
  assign _zz_4301 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_19_real));
  assign _zz_4302 = fixTo_147_dout;
  assign _zz_4303 = _zz_4304;
  assign _zz_4304 = ($signed(_zz_4305) >>> _zz_295);
  assign _zz_4305 = _zz_4306;
  assign _zz_4306 = ($signed(data_mid_17_real) - $signed(_zz_293));
  assign _zz_4307 = _zz_4308;
  assign _zz_4308 = ($signed(_zz_4309) >>> _zz_295);
  assign _zz_4309 = _zz_4310;
  assign _zz_4310 = ($signed(data_mid_17_imag) - $signed(_zz_294));
  assign _zz_4311 = _zz_4312;
  assign _zz_4312 = ($signed(_zz_4313) >>> _zz_296);
  assign _zz_4313 = _zz_4314;
  assign _zz_4314 = ($signed(data_mid_17_real) + $signed(_zz_293));
  assign _zz_4315 = _zz_4316;
  assign _zz_4316 = ($signed(_zz_4317) >>> _zz_296);
  assign _zz_4317 = _zz_4318;
  assign _zz_4318 = ($signed(data_mid_17_imag) + $signed(_zz_294));
  assign _zz_4319 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_22_real));
  assign _zz_4320 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_22_imag));
  assign _zz_4321 = fixTo_148_dout;
  assign _zz_4322 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_22_imag));
  assign _zz_4323 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_22_real));
  assign _zz_4324 = fixTo_149_dout;
  assign _zz_4325 = _zz_4326;
  assign _zz_4326 = ($signed(_zz_4327) >>> _zz_299);
  assign _zz_4327 = _zz_4328;
  assign _zz_4328 = ($signed(data_mid_20_real) - $signed(_zz_297));
  assign _zz_4329 = _zz_4330;
  assign _zz_4330 = ($signed(_zz_4331) >>> _zz_299);
  assign _zz_4331 = _zz_4332;
  assign _zz_4332 = ($signed(data_mid_20_imag) - $signed(_zz_298));
  assign _zz_4333 = _zz_4334;
  assign _zz_4334 = ($signed(_zz_4335) >>> _zz_300);
  assign _zz_4335 = _zz_4336;
  assign _zz_4336 = ($signed(data_mid_20_real) + $signed(_zz_297));
  assign _zz_4337 = _zz_4338;
  assign _zz_4338 = ($signed(_zz_4339) >>> _zz_300);
  assign _zz_4339 = _zz_4340;
  assign _zz_4340 = ($signed(data_mid_20_imag) + $signed(_zz_298));
  assign _zz_4341 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_23_real));
  assign _zz_4342 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_23_imag));
  assign _zz_4343 = fixTo_150_dout;
  assign _zz_4344 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_23_imag));
  assign _zz_4345 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_23_real));
  assign _zz_4346 = fixTo_151_dout;
  assign _zz_4347 = _zz_4348;
  assign _zz_4348 = ($signed(_zz_4349) >>> _zz_303);
  assign _zz_4349 = _zz_4350;
  assign _zz_4350 = ($signed(data_mid_21_real) - $signed(_zz_301));
  assign _zz_4351 = _zz_4352;
  assign _zz_4352 = ($signed(_zz_4353) >>> _zz_303);
  assign _zz_4353 = _zz_4354;
  assign _zz_4354 = ($signed(data_mid_21_imag) - $signed(_zz_302));
  assign _zz_4355 = _zz_4356;
  assign _zz_4356 = ($signed(_zz_4357) >>> _zz_304);
  assign _zz_4357 = _zz_4358;
  assign _zz_4358 = ($signed(data_mid_21_real) + $signed(_zz_301));
  assign _zz_4359 = _zz_4360;
  assign _zz_4360 = ($signed(_zz_4361) >>> _zz_304);
  assign _zz_4361 = _zz_4362;
  assign _zz_4362 = ($signed(data_mid_21_imag) + $signed(_zz_302));
  assign _zz_4363 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_26_real));
  assign _zz_4364 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_26_imag));
  assign _zz_4365 = fixTo_152_dout;
  assign _zz_4366 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_26_imag));
  assign _zz_4367 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_26_real));
  assign _zz_4368 = fixTo_153_dout;
  assign _zz_4369 = _zz_4370;
  assign _zz_4370 = ($signed(_zz_4371) >>> _zz_307);
  assign _zz_4371 = _zz_4372;
  assign _zz_4372 = ($signed(data_mid_24_real) - $signed(_zz_305));
  assign _zz_4373 = _zz_4374;
  assign _zz_4374 = ($signed(_zz_4375) >>> _zz_307);
  assign _zz_4375 = _zz_4376;
  assign _zz_4376 = ($signed(data_mid_24_imag) - $signed(_zz_306));
  assign _zz_4377 = _zz_4378;
  assign _zz_4378 = ($signed(_zz_4379) >>> _zz_308);
  assign _zz_4379 = _zz_4380;
  assign _zz_4380 = ($signed(data_mid_24_real) + $signed(_zz_305));
  assign _zz_4381 = _zz_4382;
  assign _zz_4382 = ($signed(_zz_4383) >>> _zz_308);
  assign _zz_4383 = _zz_4384;
  assign _zz_4384 = ($signed(data_mid_24_imag) + $signed(_zz_306));
  assign _zz_4385 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_27_real));
  assign _zz_4386 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_27_imag));
  assign _zz_4387 = fixTo_154_dout;
  assign _zz_4388 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_27_imag));
  assign _zz_4389 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_27_real));
  assign _zz_4390 = fixTo_155_dout;
  assign _zz_4391 = _zz_4392;
  assign _zz_4392 = ($signed(_zz_4393) >>> _zz_311);
  assign _zz_4393 = _zz_4394;
  assign _zz_4394 = ($signed(data_mid_25_real) - $signed(_zz_309));
  assign _zz_4395 = _zz_4396;
  assign _zz_4396 = ($signed(_zz_4397) >>> _zz_311);
  assign _zz_4397 = _zz_4398;
  assign _zz_4398 = ($signed(data_mid_25_imag) - $signed(_zz_310));
  assign _zz_4399 = _zz_4400;
  assign _zz_4400 = ($signed(_zz_4401) >>> _zz_312);
  assign _zz_4401 = _zz_4402;
  assign _zz_4402 = ($signed(data_mid_25_real) + $signed(_zz_309));
  assign _zz_4403 = _zz_4404;
  assign _zz_4404 = ($signed(_zz_4405) >>> _zz_312);
  assign _zz_4405 = _zz_4406;
  assign _zz_4406 = ($signed(data_mid_25_imag) + $signed(_zz_310));
  assign _zz_4407 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_30_real));
  assign _zz_4408 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_30_imag));
  assign _zz_4409 = fixTo_156_dout;
  assign _zz_4410 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_30_imag));
  assign _zz_4411 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_30_real));
  assign _zz_4412 = fixTo_157_dout;
  assign _zz_4413 = _zz_4414;
  assign _zz_4414 = ($signed(_zz_4415) >>> _zz_315);
  assign _zz_4415 = _zz_4416;
  assign _zz_4416 = ($signed(data_mid_28_real) - $signed(_zz_313));
  assign _zz_4417 = _zz_4418;
  assign _zz_4418 = ($signed(_zz_4419) >>> _zz_315);
  assign _zz_4419 = _zz_4420;
  assign _zz_4420 = ($signed(data_mid_28_imag) - $signed(_zz_314));
  assign _zz_4421 = _zz_4422;
  assign _zz_4422 = ($signed(_zz_4423) >>> _zz_316);
  assign _zz_4423 = _zz_4424;
  assign _zz_4424 = ($signed(data_mid_28_real) + $signed(_zz_313));
  assign _zz_4425 = _zz_4426;
  assign _zz_4426 = ($signed(_zz_4427) >>> _zz_316);
  assign _zz_4427 = _zz_4428;
  assign _zz_4428 = ($signed(data_mid_28_imag) + $signed(_zz_314));
  assign _zz_4429 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_31_real));
  assign _zz_4430 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_31_imag));
  assign _zz_4431 = fixTo_158_dout;
  assign _zz_4432 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_31_imag));
  assign _zz_4433 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_31_real));
  assign _zz_4434 = fixTo_159_dout;
  assign _zz_4435 = _zz_4436;
  assign _zz_4436 = ($signed(_zz_4437) >>> _zz_319);
  assign _zz_4437 = _zz_4438;
  assign _zz_4438 = ($signed(data_mid_29_real) - $signed(_zz_317));
  assign _zz_4439 = _zz_4440;
  assign _zz_4440 = ($signed(_zz_4441) >>> _zz_319);
  assign _zz_4441 = _zz_4442;
  assign _zz_4442 = ($signed(data_mid_29_imag) - $signed(_zz_318));
  assign _zz_4443 = _zz_4444;
  assign _zz_4444 = ($signed(_zz_4445) >>> _zz_320);
  assign _zz_4445 = _zz_4446;
  assign _zz_4446 = ($signed(data_mid_29_real) + $signed(_zz_317));
  assign _zz_4447 = _zz_4448;
  assign _zz_4448 = ($signed(_zz_4449) >>> _zz_320);
  assign _zz_4449 = _zz_4450;
  assign _zz_4450 = ($signed(data_mid_29_imag) + $signed(_zz_318));
  assign _zz_4451 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_34_real));
  assign _zz_4452 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_34_imag));
  assign _zz_4453 = fixTo_160_dout;
  assign _zz_4454 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_34_imag));
  assign _zz_4455 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_34_real));
  assign _zz_4456 = fixTo_161_dout;
  assign _zz_4457 = _zz_4458;
  assign _zz_4458 = ($signed(_zz_4459) >>> _zz_323);
  assign _zz_4459 = _zz_4460;
  assign _zz_4460 = ($signed(data_mid_32_real) - $signed(_zz_321));
  assign _zz_4461 = _zz_4462;
  assign _zz_4462 = ($signed(_zz_4463) >>> _zz_323);
  assign _zz_4463 = _zz_4464;
  assign _zz_4464 = ($signed(data_mid_32_imag) - $signed(_zz_322));
  assign _zz_4465 = _zz_4466;
  assign _zz_4466 = ($signed(_zz_4467) >>> _zz_324);
  assign _zz_4467 = _zz_4468;
  assign _zz_4468 = ($signed(data_mid_32_real) + $signed(_zz_321));
  assign _zz_4469 = _zz_4470;
  assign _zz_4470 = ($signed(_zz_4471) >>> _zz_324);
  assign _zz_4471 = _zz_4472;
  assign _zz_4472 = ($signed(data_mid_32_imag) + $signed(_zz_322));
  assign _zz_4473 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_35_real));
  assign _zz_4474 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_35_imag));
  assign _zz_4475 = fixTo_162_dout;
  assign _zz_4476 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_35_imag));
  assign _zz_4477 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_35_real));
  assign _zz_4478 = fixTo_163_dout;
  assign _zz_4479 = _zz_4480;
  assign _zz_4480 = ($signed(_zz_4481) >>> _zz_327);
  assign _zz_4481 = _zz_4482;
  assign _zz_4482 = ($signed(data_mid_33_real) - $signed(_zz_325));
  assign _zz_4483 = _zz_4484;
  assign _zz_4484 = ($signed(_zz_4485) >>> _zz_327);
  assign _zz_4485 = _zz_4486;
  assign _zz_4486 = ($signed(data_mid_33_imag) - $signed(_zz_326));
  assign _zz_4487 = _zz_4488;
  assign _zz_4488 = ($signed(_zz_4489) >>> _zz_328);
  assign _zz_4489 = _zz_4490;
  assign _zz_4490 = ($signed(data_mid_33_real) + $signed(_zz_325));
  assign _zz_4491 = _zz_4492;
  assign _zz_4492 = ($signed(_zz_4493) >>> _zz_328);
  assign _zz_4493 = _zz_4494;
  assign _zz_4494 = ($signed(data_mid_33_imag) + $signed(_zz_326));
  assign _zz_4495 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_38_real));
  assign _zz_4496 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_38_imag));
  assign _zz_4497 = fixTo_164_dout;
  assign _zz_4498 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_38_imag));
  assign _zz_4499 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_38_real));
  assign _zz_4500 = fixTo_165_dout;
  assign _zz_4501 = _zz_4502;
  assign _zz_4502 = ($signed(_zz_4503) >>> _zz_331);
  assign _zz_4503 = _zz_4504;
  assign _zz_4504 = ($signed(data_mid_36_real) - $signed(_zz_329));
  assign _zz_4505 = _zz_4506;
  assign _zz_4506 = ($signed(_zz_4507) >>> _zz_331);
  assign _zz_4507 = _zz_4508;
  assign _zz_4508 = ($signed(data_mid_36_imag) - $signed(_zz_330));
  assign _zz_4509 = _zz_4510;
  assign _zz_4510 = ($signed(_zz_4511) >>> _zz_332);
  assign _zz_4511 = _zz_4512;
  assign _zz_4512 = ($signed(data_mid_36_real) + $signed(_zz_329));
  assign _zz_4513 = _zz_4514;
  assign _zz_4514 = ($signed(_zz_4515) >>> _zz_332);
  assign _zz_4515 = _zz_4516;
  assign _zz_4516 = ($signed(data_mid_36_imag) + $signed(_zz_330));
  assign _zz_4517 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_39_real));
  assign _zz_4518 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_39_imag));
  assign _zz_4519 = fixTo_166_dout;
  assign _zz_4520 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_39_imag));
  assign _zz_4521 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_39_real));
  assign _zz_4522 = fixTo_167_dout;
  assign _zz_4523 = _zz_4524;
  assign _zz_4524 = ($signed(_zz_4525) >>> _zz_335);
  assign _zz_4525 = _zz_4526;
  assign _zz_4526 = ($signed(data_mid_37_real) - $signed(_zz_333));
  assign _zz_4527 = _zz_4528;
  assign _zz_4528 = ($signed(_zz_4529) >>> _zz_335);
  assign _zz_4529 = _zz_4530;
  assign _zz_4530 = ($signed(data_mid_37_imag) - $signed(_zz_334));
  assign _zz_4531 = _zz_4532;
  assign _zz_4532 = ($signed(_zz_4533) >>> _zz_336);
  assign _zz_4533 = _zz_4534;
  assign _zz_4534 = ($signed(data_mid_37_real) + $signed(_zz_333));
  assign _zz_4535 = _zz_4536;
  assign _zz_4536 = ($signed(_zz_4537) >>> _zz_336);
  assign _zz_4537 = _zz_4538;
  assign _zz_4538 = ($signed(data_mid_37_imag) + $signed(_zz_334));
  assign _zz_4539 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_42_real));
  assign _zz_4540 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_42_imag));
  assign _zz_4541 = fixTo_168_dout;
  assign _zz_4542 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_42_imag));
  assign _zz_4543 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_42_real));
  assign _zz_4544 = fixTo_169_dout;
  assign _zz_4545 = _zz_4546;
  assign _zz_4546 = ($signed(_zz_4547) >>> _zz_339);
  assign _zz_4547 = _zz_4548;
  assign _zz_4548 = ($signed(data_mid_40_real) - $signed(_zz_337));
  assign _zz_4549 = _zz_4550;
  assign _zz_4550 = ($signed(_zz_4551) >>> _zz_339);
  assign _zz_4551 = _zz_4552;
  assign _zz_4552 = ($signed(data_mid_40_imag) - $signed(_zz_338));
  assign _zz_4553 = _zz_4554;
  assign _zz_4554 = ($signed(_zz_4555) >>> _zz_340);
  assign _zz_4555 = _zz_4556;
  assign _zz_4556 = ($signed(data_mid_40_real) + $signed(_zz_337));
  assign _zz_4557 = _zz_4558;
  assign _zz_4558 = ($signed(_zz_4559) >>> _zz_340);
  assign _zz_4559 = _zz_4560;
  assign _zz_4560 = ($signed(data_mid_40_imag) + $signed(_zz_338));
  assign _zz_4561 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_43_real));
  assign _zz_4562 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_43_imag));
  assign _zz_4563 = fixTo_170_dout;
  assign _zz_4564 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_43_imag));
  assign _zz_4565 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_43_real));
  assign _zz_4566 = fixTo_171_dout;
  assign _zz_4567 = _zz_4568;
  assign _zz_4568 = ($signed(_zz_4569) >>> _zz_343);
  assign _zz_4569 = _zz_4570;
  assign _zz_4570 = ($signed(data_mid_41_real) - $signed(_zz_341));
  assign _zz_4571 = _zz_4572;
  assign _zz_4572 = ($signed(_zz_4573) >>> _zz_343);
  assign _zz_4573 = _zz_4574;
  assign _zz_4574 = ($signed(data_mid_41_imag) - $signed(_zz_342));
  assign _zz_4575 = _zz_4576;
  assign _zz_4576 = ($signed(_zz_4577) >>> _zz_344);
  assign _zz_4577 = _zz_4578;
  assign _zz_4578 = ($signed(data_mid_41_real) + $signed(_zz_341));
  assign _zz_4579 = _zz_4580;
  assign _zz_4580 = ($signed(_zz_4581) >>> _zz_344);
  assign _zz_4581 = _zz_4582;
  assign _zz_4582 = ($signed(data_mid_41_imag) + $signed(_zz_342));
  assign _zz_4583 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_46_real));
  assign _zz_4584 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_46_imag));
  assign _zz_4585 = fixTo_172_dout;
  assign _zz_4586 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_46_imag));
  assign _zz_4587 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_46_real));
  assign _zz_4588 = fixTo_173_dout;
  assign _zz_4589 = _zz_4590;
  assign _zz_4590 = ($signed(_zz_4591) >>> _zz_347);
  assign _zz_4591 = _zz_4592;
  assign _zz_4592 = ($signed(data_mid_44_real) - $signed(_zz_345));
  assign _zz_4593 = _zz_4594;
  assign _zz_4594 = ($signed(_zz_4595) >>> _zz_347);
  assign _zz_4595 = _zz_4596;
  assign _zz_4596 = ($signed(data_mid_44_imag) - $signed(_zz_346));
  assign _zz_4597 = _zz_4598;
  assign _zz_4598 = ($signed(_zz_4599) >>> _zz_348);
  assign _zz_4599 = _zz_4600;
  assign _zz_4600 = ($signed(data_mid_44_real) + $signed(_zz_345));
  assign _zz_4601 = _zz_4602;
  assign _zz_4602 = ($signed(_zz_4603) >>> _zz_348);
  assign _zz_4603 = _zz_4604;
  assign _zz_4604 = ($signed(data_mid_44_imag) + $signed(_zz_346));
  assign _zz_4605 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_47_real));
  assign _zz_4606 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_47_imag));
  assign _zz_4607 = fixTo_174_dout;
  assign _zz_4608 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_47_imag));
  assign _zz_4609 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_47_real));
  assign _zz_4610 = fixTo_175_dout;
  assign _zz_4611 = _zz_4612;
  assign _zz_4612 = ($signed(_zz_4613) >>> _zz_351);
  assign _zz_4613 = _zz_4614;
  assign _zz_4614 = ($signed(data_mid_45_real) - $signed(_zz_349));
  assign _zz_4615 = _zz_4616;
  assign _zz_4616 = ($signed(_zz_4617) >>> _zz_351);
  assign _zz_4617 = _zz_4618;
  assign _zz_4618 = ($signed(data_mid_45_imag) - $signed(_zz_350));
  assign _zz_4619 = _zz_4620;
  assign _zz_4620 = ($signed(_zz_4621) >>> _zz_352);
  assign _zz_4621 = _zz_4622;
  assign _zz_4622 = ($signed(data_mid_45_real) + $signed(_zz_349));
  assign _zz_4623 = _zz_4624;
  assign _zz_4624 = ($signed(_zz_4625) >>> _zz_352);
  assign _zz_4625 = _zz_4626;
  assign _zz_4626 = ($signed(data_mid_45_imag) + $signed(_zz_350));
  assign _zz_4627 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_50_real));
  assign _zz_4628 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_50_imag));
  assign _zz_4629 = fixTo_176_dout;
  assign _zz_4630 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_50_imag));
  assign _zz_4631 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_50_real));
  assign _zz_4632 = fixTo_177_dout;
  assign _zz_4633 = _zz_4634;
  assign _zz_4634 = ($signed(_zz_4635) >>> _zz_355);
  assign _zz_4635 = _zz_4636;
  assign _zz_4636 = ($signed(data_mid_48_real) - $signed(_zz_353));
  assign _zz_4637 = _zz_4638;
  assign _zz_4638 = ($signed(_zz_4639) >>> _zz_355);
  assign _zz_4639 = _zz_4640;
  assign _zz_4640 = ($signed(data_mid_48_imag) - $signed(_zz_354));
  assign _zz_4641 = _zz_4642;
  assign _zz_4642 = ($signed(_zz_4643) >>> _zz_356);
  assign _zz_4643 = _zz_4644;
  assign _zz_4644 = ($signed(data_mid_48_real) + $signed(_zz_353));
  assign _zz_4645 = _zz_4646;
  assign _zz_4646 = ($signed(_zz_4647) >>> _zz_356);
  assign _zz_4647 = _zz_4648;
  assign _zz_4648 = ($signed(data_mid_48_imag) + $signed(_zz_354));
  assign _zz_4649 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_51_real));
  assign _zz_4650 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_51_imag));
  assign _zz_4651 = fixTo_178_dout;
  assign _zz_4652 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_51_imag));
  assign _zz_4653 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_51_real));
  assign _zz_4654 = fixTo_179_dout;
  assign _zz_4655 = _zz_4656;
  assign _zz_4656 = ($signed(_zz_4657) >>> _zz_359);
  assign _zz_4657 = _zz_4658;
  assign _zz_4658 = ($signed(data_mid_49_real) - $signed(_zz_357));
  assign _zz_4659 = _zz_4660;
  assign _zz_4660 = ($signed(_zz_4661) >>> _zz_359);
  assign _zz_4661 = _zz_4662;
  assign _zz_4662 = ($signed(data_mid_49_imag) - $signed(_zz_358));
  assign _zz_4663 = _zz_4664;
  assign _zz_4664 = ($signed(_zz_4665) >>> _zz_360);
  assign _zz_4665 = _zz_4666;
  assign _zz_4666 = ($signed(data_mid_49_real) + $signed(_zz_357));
  assign _zz_4667 = _zz_4668;
  assign _zz_4668 = ($signed(_zz_4669) >>> _zz_360);
  assign _zz_4669 = _zz_4670;
  assign _zz_4670 = ($signed(data_mid_49_imag) + $signed(_zz_358));
  assign _zz_4671 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_54_real));
  assign _zz_4672 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_54_imag));
  assign _zz_4673 = fixTo_180_dout;
  assign _zz_4674 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_54_imag));
  assign _zz_4675 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_54_real));
  assign _zz_4676 = fixTo_181_dout;
  assign _zz_4677 = _zz_4678;
  assign _zz_4678 = ($signed(_zz_4679) >>> _zz_363);
  assign _zz_4679 = _zz_4680;
  assign _zz_4680 = ($signed(data_mid_52_real) - $signed(_zz_361));
  assign _zz_4681 = _zz_4682;
  assign _zz_4682 = ($signed(_zz_4683) >>> _zz_363);
  assign _zz_4683 = _zz_4684;
  assign _zz_4684 = ($signed(data_mid_52_imag) - $signed(_zz_362));
  assign _zz_4685 = _zz_4686;
  assign _zz_4686 = ($signed(_zz_4687) >>> _zz_364);
  assign _zz_4687 = _zz_4688;
  assign _zz_4688 = ($signed(data_mid_52_real) + $signed(_zz_361));
  assign _zz_4689 = _zz_4690;
  assign _zz_4690 = ($signed(_zz_4691) >>> _zz_364);
  assign _zz_4691 = _zz_4692;
  assign _zz_4692 = ($signed(data_mid_52_imag) + $signed(_zz_362));
  assign _zz_4693 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_55_real));
  assign _zz_4694 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_55_imag));
  assign _zz_4695 = fixTo_182_dout;
  assign _zz_4696 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_55_imag));
  assign _zz_4697 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_55_real));
  assign _zz_4698 = fixTo_183_dout;
  assign _zz_4699 = _zz_4700;
  assign _zz_4700 = ($signed(_zz_4701) >>> _zz_367);
  assign _zz_4701 = _zz_4702;
  assign _zz_4702 = ($signed(data_mid_53_real) - $signed(_zz_365));
  assign _zz_4703 = _zz_4704;
  assign _zz_4704 = ($signed(_zz_4705) >>> _zz_367);
  assign _zz_4705 = _zz_4706;
  assign _zz_4706 = ($signed(data_mid_53_imag) - $signed(_zz_366));
  assign _zz_4707 = _zz_4708;
  assign _zz_4708 = ($signed(_zz_4709) >>> _zz_368);
  assign _zz_4709 = _zz_4710;
  assign _zz_4710 = ($signed(data_mid_53_real) + $signed(_zz_365));
  assign _zz_4711 = _zz_4712;
  assign _zz_4712 = ($signed(_zz_4713) >>> _zz_368);
  assign _zz_4713 = _zz_4714;
  assign _zz_4714 = ($signed(data_mid_53_imag) + $signed(_zz_366));
  assign _zz_4715 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_58_real));
  assign _zz_4716 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_58_imag));
  assign _zz_4717 = fixTo_184_dout;
  assign _zz_4718 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_58_imag));
  assign _zz_4719 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_58_real));
  assign _zz_4720 = fixTo_185_dout;
  assign _zz_4721 = _zz_4722;
  assign _zz_4722 = ($signed(_zz_4723) >>> _zz_371);
  assign _zz_4723 = _zz_4724;
  assign _zz_4724 = ($signed(data_mid_56_real) - $signed(_zz_369));
  assign _zz_4725 = _zz_4726;
  assign _zz_4726 = ($signed(_zz_4727) >>> _zz_371);
  assign _zz_4727 = _zz_4728;
  assign _zz_4728 = ($signed(data_mid_56_imag) - $signed(_zz_370));
  assign _zz_4729 = _zz_4730;
  assign _zz_4730 = ($signed(_zz_4731) >>> _zz_372);
  assign _zz_4731 = _zz_4732;
  assign _zz_4732 = ($signed(data_mid_56_real) + $signed(_zz_369));
  assign _zz_4733 = _zz_4734;
  assign _zz_4734 = ($signed(_zz_4735) >>> _zz_372);
  assign _zz_4735 = _zz_4736;
  assign _zz_4736 = ($signed(data_mid_56_imag) + $signed(_zz_370));
  assign _zz_4737 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_59_real));
  assign _zz_4738 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_59_imag));
  assign _zz_4739 = fixTo_186_dout;
  assign _zz_4740 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_59_imag));
  assign _zz_4741 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_59_real));
  assign _zz_4742 = fixTo_187_dout;
  assign _zz_4743 = _zz_4744;
  assign _zz_4744 = ($signed(_zz_4745) >>> _zz_375);
  assign _zz_4745 = _zz_4746;
  assign _zz_4746 = ($signed(data_mid_57_real) - $signed(_zz_373));
  assign _zz_4747 = _zz_4748;
  assign _zz_4748 = ($signed(_zz_4749) >>> _zz_375);
  assign _zz_4749 = _zz_4750;
  assign _zz_4750 = ($signed(data_mid_57_imag) - $signed(_zz_374));
  assign _zz_4751 = _zz_4752;
  assign _zz_4752 = ($signed(_zz_4753) >>> _zz_376);
  assign _zz_4753 = _zz_4754;
  assign _zz_4754 = ($signed(data_mid_57_real) + $signed(_zz_373));
  assign _zz_4755 = _zz_4756;
  assign _zz_4756 = ($signed(_zz_4757) >>> _zz_376);
  assign _zz_4757 = _zz_4758;
  assign _zz_4758 = ($signed(data_mid_57_imag) + $signed(_zz_374));
  assign _zz_4759 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_62_real));
  assign _zz_4760 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_62_imag));
  assign _zz_4761 = fixTo_188_dout;
  assign _zz_4762 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_62_imag));
  assign _zz_4763 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_62_real));
  assign _zz_4764 = fixTo_189_dout;
  assign _zz_4765 = _zz_4766;
  assign _zz_4766 = ($signed(_zz_4767) >>> _zz_379);
  assign _zz_4767 = _zz_4768;
  assign _zz_4768 = ($signed(data_mid_60_real) - $signed(_zz_377));
  assign _zz_4769 = _zz_4770;
  assign _zz_4770 = ($signed(_zz_4771) >>> _zz_379);
  assign _zz_4771 = _zz_4772;
  assign _zz_4772 = ($signed(data_mid_60_imag) - $signed(_zz_378));
  assign _zz_4773 = _zz_4774;
  assign _zz_4774 = ($signed(_zz_4775) >>> _zz_380);
  assign _zz_4775 = _zz_4776;
  assign _zz_4776 = ($signed(data_mid_60_real) + $signed(_zz_377));
  assign _zz_4777 = _zz_4778;
  assign _zz_4778 = ($signed(_zz_4779) >>> _zz_380);
  assign _zz_4779 = _zz_4780;
  assign _zz_4780 = ($signed(data_mid_60_imag) + $signed(_zz_378));
  assign _zz_4781 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_63_real));
  assign _zz_4782 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_63_imag));
  assign _zz_4783 = fixTo_190_dout;
  assign _zz_4784 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_63_imag));
  assign _zz_4785 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_63_real));
  assign _zz_4786 = fixTo_191_dout;
  assign _zz_4787 = _zz_4788;
  assign _zz_4788 = ($signed(_zz_4789) >>> _zz_383);
  assign _zz_4789 = _zz_4790;
  assign _zz_4790 = ($signed(data_mid_61_real) - $signed(_zz_381));
  assign _zz_4791 = _zz_4792;
  assign _zz_4792 = ($signed(_zz_4793) >>> _zz_383);
  assign _zz_4793 = _zz_4794;
  assign _zz_4794 = ($signed(data_mid_61_imag) - $signed(_zz_382));
  assign _zz_4795 = _zz_4796;
  assign _zz_4796 = ($signed(_zz_4797) >>> _zz_384);
  assign _zz_4797 = _zz_4798;
  assign _zz_4798 = ($signed(data_mid_61_real) + $signed(_zz_381));
  assign _zz_4799 = _zz_4800;
  assign _zz_4800 = ($signed(_zz_4801) >>> _zz_384);
  assign _zz_4801 = _zz_4802;
  assign _zz_4802 = ($signed(data_mid_61_imag) + $signed(_zz_382));
  assign _zz_4803 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_66_real));
  assign _zz_4804 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_66_imag));
  assign _zz_4805 = fixTo_192_dout;
  assign _zz_4806 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_66_imag));
  assign _zz_4807 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_66_real));
  assign _zz_4808 = fixTo_193_dout;
  assign _zz_4809 = _zz_4810;
  assign _zz_4810 = ($signed(_zz_4811) >>> _zz_387);
  assign _zz_4811 = _zz_4812;
  assign _zz_4812 = ($signed(data_mid_64_real) - $signed(_zz_385));
  assign _zz_4813 = _zz_4814;
  assign _zz_4814 = ($signed(_zz_4815) >>> _zz_387);
  assign _zz_4815 = _zz_4816;
  assign _zz_4816 = ($signed(data_mid_64_imag) - $signed(_zz_386));
  assign _zz_4817 = _zz_4818;
  assign _zz_4818 = ($signed(_zz_4819) >>> _zz_388);
  assign _zz_4819 = _zz_4820;
  assign _zz_4820 = ($signed(data_mid_64_real) + $signed(_zz_385));
  assign _zz_4821 = _zz_4822;
  assign _zz_4822 = ($signed(_zz_4823) >>> _zz_388);
  assign _zz_4823 = _zz_4824;
  assign _zz_4824 = ($signed(data_mid_64_imag) + $signed(_zz_386));
  assign _zz_4825 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_67_real));
  assign _zz_4826 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_67_imag));
  assign _zz_4827 = fixTo_194_dout;
  assign _zz_4828 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_67_imag));
  assign _zz_4829 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_67_real));
  assign _zz_4830 = fixTo_195_dout;
  assign _zz_4831 = _zz_4832;
  assign _zz_4832 = ($signed(_zz_4833) >>> _zz_391);
  assign _zz_4833 = _zz_4834;
  assign _zz_4834 = ($signed(data_mid_65_real) - $signed(_zz_389));
  assign _zz_4835 = _zz_4836;
  assign _zz_4836 = ($signed(_zz_4837) >>> _zz_391);
  assign _zz_4837 = _zz_4838;
  assign _zz_4838 = ($signed(data_mid_65_imag) - $signed(_zz_390));
  assign _zz_4839 = _zz_4840;
  assign _zz_4840 = ($signed(_zz_4841) >>> _zz_392);
  assign _zz_4841 = _zz_4842;
  assign _zz_4842 = ($signed(data_mid_65_real) + $signed(_zz_389));
  assign _zz_4843 = _zz_4844;
  assign _zz_4844 = ($signed(_zz_4845) >>> _zz_392);
  assign _zz_4845 = _zz_4846;
  assign _zz_4846 = ($signed(data_mid_65_imag) + $signed(_zz_390));
  assign _zz_4847 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_70_real));
  assign _zz_4848 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_70_imag));
  assign _zz_4849 = fixTo_196_dout;
  assign _zz_4850 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_70_imag));
  assign _zz_4851 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_70_real));
  assign _zz_4852 = fixTo_197_dout;
  assign _zz_4853 = _zz_4854;
  assign _zz_4854 = ($signed(_zz_4855) >>> _zz_395);
  assign _zz_4855 = _zz_4856;
  assign _zz_4856 = ($signed(data_mid_68_real) - $signed(_zz_393));
  assign _zz_4857 = _zz_4858;
  assign _zz_4858 = ($signed(_zz_4859) >>> _zz_395);
  assign _zz_4859 = _zz_4860;
  assign _zz_4860 = ($signed(data_mid_68_imag) - $signed(_zz_394));
  assign _zz_4861 = _zz_4862;
  assign _zz_4862 = ($signed(_zz_4863) >>> _zz_396);
  assign _zz_4863 = _zz_4864;
  assign _zz_4864 = ($signed(data_mid_68_real) + $signed(_zz_393));
  assign _zz_4865 = _zz_4866;
  assign _zz_4866 = ($signed(_zz_4867) >>> _zz_396);
  assign _zz_4867 = _zz_4868;
  assign _zz_4868 = ($signed(data_mid_68_imag) + $signed(_zz_394));
  assign _zz_4869 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_71_real));
  assign _zz_4870 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_71_imag));
  assign _zz_4871 = fixTo_198_dout;
  assign _zz_4872 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_71_imag));
  assign _zz_4873 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_71_real));
  assign _zz_4874 = fixTo_199_dout;
  assign _zz_4875 = _zz_4876;
  assign _zz_4876 = ($signed(_zz_4877) >>> _zz_399);
  assign _zz_4877 = _zz_4878;
  assign _zz_4878 = ($signed(data_mid_69_real) - $signed(_zz_397));
  assign _zz_4879 = _zz_4880;
  assign _zz_4880 = ($signed(_zz_4881) >>> _zz_399);
  assign _zz_4881 = _zz_4882;
  assign _zz_4882 = ($signed(data_mid_69_imag) - $signed(_zz_398));
  assign _zz_4883 = _zz_4884;
  assign _zz_4884 = ($signed(_zz_4885) >>> _zz_400);
  assign _zz_4885 = _zz_4886;
  assign _zz_4886 = ($signed(data_mid_69_real) + $signed(_zz_397));
  assign _zz_4887 = _zz_4888;
  assign _zz_4888 = ($signed(_zz_4889) >>> _zz_400);
  assign _zz_4889 = _zz_4890;
  assign _zz_4890 = ($signed(data_mid_69_imag) + $signed(_zz_398));
  assign _zz_4891 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_74_real));
  assign _zz_4892 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_74_imag));
  assign _zz_4893 = fixTo_200_dout;
  assign _zz_4894 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_74_imag));
  assign _zz_4895 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_74_real));
  assign _zz_4896 = fixTo_201_dout;
  assign _zz_4897 = _zz_4898;
  assign _zz_4898 = ($signed(_zz_4899) >>> _zz_403);
  assign _zz_4899 = _zz_4900;
  assign _zz_4900 = ($signed(data_mid_72_real) - $signed(_zz_401));
  assign _zz_4901 = _zz_4902;
  assign _zz_4902 = ($signed(_zz_4903) >>> _zz_403);
  assign _zz_4903 = _zz_4904;
  assign _zz_4904 = ($signed(data_mid_72_imag) - $signed(_zz_402));
  assign _zz_4905 = _zz_4906;
  assign _zz_4906 = ($signed(_zz_4907) >>> _zz_404);
  assign _zz_4907 = _zz_4908;
  assign _zz_4908 = ($signed(data_mid_72_real) + $signed(_zz_401));
  assign _zz_4909 = _zz_4910;
  assign _zz_4910 = ($signed(_zz_4911) >>> _zz_404);
  assign _zz_4911 = _zz_4912;
  assign _zz_4912 = ($signed(data_mid_72_imag) + $signed(_zz_402));
  assign _zz_4913 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_75_real));
  assign _zz_4914 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_75_imag));
  assign _zz_4915 = fixTo_202_dout;
  assign _zz_4916 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_75_imag));
  assign _zz_4917 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_75_real));
  assign _zz_4918 = fixTo_203_dout;
  assign _zz_4919 = _zz_4920;
  assign _zz_4920 = ($signed(_zz_4921) >>> _zz_407);
  assign _zz_4921 = _zz_4922;
  assign _zz_4922 = ($signed(data_mid_73_real) - $signed(_zz_405));
  assign _zz_4923 = _zz_4924;
  assign _zz_4924 = ($signed(_zz_4925) >>> _zz_407);
  assign _zz_4925 = _zz_4926;
  assign _zz_4926 = ($signed(data_mid_73_imag) - $signed(_zz_406));
  assign _zz_4927 = _zz_4928;
  assign _zz_4928 = ($signed(_zz_4929) >>> _zz_408);
  assign _zz_4929 = _zz_4930;
  assign _zz_4930 = ($signed(data_mid_73_real) + $signed(_zz_405));
  assign _zz_4931 = _zz_4932;
  assign _zz_4932 = ($signed(_zz_4933) >>> _zz_408);
  assign _zz_4933 = _zz_4934;
  assign _zz_4934 = ($signed(data_mid_73_imag) + $signed(_zz_406));
  assign _zz_4935 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_78_real));
  assign _zz_4936 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_78_imag));
  assign _zz_4937 = fixTo_204_dout;
  assign _zz_4938 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_78_imag));
  assign _zz_4939 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_78_real));
  assign _zz_4940 = fixTo_205_dout;
  assign _zz_4941 = _zz_4942;
  assign _zz_4942 = ($signed(_zz_4943) >>> _zz_411);
  assign _zz_4943 = _zz_4944;
  assign _zz_4944 = ($signed(data_mid_76_real) - $signed(_zz_409));
  assign _zz_4945 = _zz_4946;
  assign _zz_4946 = ($signed(_zz_4947) >>> _zz_411);
  assign _zz_4947 = _zz_4948;
  assign _zz_4948 = ($signed(data_mid_76_imag) - $signed(_zz_410));
  assign _zz_4949 = _zz_4950;
  assign _zz_4950 = ($signed(_zz_4951) >>> _zz_412);
  assign _zz_4951 = _zz_4952;
  assign _zz_4952 = ($signed(data_mid_76_real) + $signed(_zz_409));
  assign _zz_4953 = _zz_4954;
  assign _zz_4954 = ($signed(_zz_4955) >>> _zz_412);
  assign _zz_4955 = _zz_4956;
  assign _zz_4956 = ($signed(data_mid_76_imag) + $signed(_zz_410));
  assign _zz_4957 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_79_real));
  assign _zz_4958 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_79_imag));
  assign _zz_4959 = fixTo_206_dout;
  assign _zz_4960 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_79_imag));
  assign _zz_4961 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_79_real));
  assign _zz_4962 = fixTo_207_dout;
  assign _zz_4963 = _zz_4964;
  assign _zz_4964 = ($signed(_zz_4965) >>> _zz_415);
  assign _zz_4965 = _zz_4966;
  assign _zz_4966 = ($signed(data_mid_77_real) - $signed(_zz_413));
  assign _zz_4967 = _zz_4968;
  assign _zz_4968 = ($signed(_zz_4969) >>> _zz_415);
  assign _zz_4969 = _zz_4970;
  assign _zz_4970 = ($signed(data_mid_77_imag) - $signed(_zz_414));
  assign _zz_4971 = _zz_4972;
  assign _zz_4972 = ($signed(_zz_4973) >>> _zz_416);
  assign _zz_4973 = _zz_4974;
  assign _zz_4974 = ($signed(data_mid_77_real) + $signed(_zz_413));
  assign _zz_4975 = _zz_4976;
  assign _zz_4976 = ($signed(_zz_4977) >>> _zz_416);
  assign _zz_4977 = _zz_4978;
  assign _zz_4978 = ($signed(data_mid_77_imag) + $signed(_zz_414));
  assign _zz_4979 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_82_real));
  assign _zz_4980 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_82_imag));
  assign _zz_4981 = fixTo_208_dout;
  assign _zz_4982 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_82_imag));
  assign _zz_4983 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_82_real));
  assign _zz_4984 = fixTo_209_dout;
  assign _zz_4985 = _zz_4986;
  assign _zz_4986 = ($signed(_zz_4987) >>> _zz_419);
  assign _zz_4987 = _zz_4988;
  assign _zz_4988 = ($signed(data_mid_80_real) - $signed(_zz_417));
  assign _zz_4989 = _zz_4990;
  assign _zz_4990 = ($signed(_zz_4991) >>> _zz_419);
  assign _zz_4991 = _zz_4992;
  assign _zz_4992 = ($signed(data_mid_80_imag) - $signed(_zz_418));
  assign _zz_4993 = _zz_4994;
  assign _zz_4994 = ($signed(_zz_4995) >>> _zz_420);
  assign _zz_4995 = _zz_4996;
  assign _zz_4996 = ($signed(data_mid_80_real) + $signed(_zz_417));
  assign _zz_4997 = _zz_4998;
  assign _zz_4998 = ($signed(_zz_4999) >>> _zz_420);
  assign _zz_4999 = _zz_5000;
  assign _zz_5000 = ($signed(data_mid_80_imag) + $signed(_zz_418));
  assign _zz_5001 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_83_real));
  assign _zz_5002 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_83_imag));
  assign _zz_5003 = fixTo_210_dout;
  assign _zz_5004 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_83_imag));
  assign _zz_5005 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_83_real));
  assign _zz_5006 = fixTo_211_dout;
  assign _zz_5007 = _zz_5008;
  assign _zz_5008 = ($signed(_zz_5009) >>> _zz_423);
  assign _zz_5009 = _zz_5010;
  assign _zz_5010 = ($signed(data_mid_81_real) - $signed(_zz_421));
  assign _zz_5011 = _zz_5012;
  assign _zz_5012 = ($signed(_zz_5013) >>> _zz_423);
  assign _zz_5013 = _zz_5014;
  assign _zz_5014 = ($signed(data_mid_81_imag) - $signed(_zz_422));
  assign _zz_5015 = _zz_5016;
  assign _zz_5016 = ($signed(_zz_5017) >>> _zz_424);
  assign _zz_5017 = _zz_5018;
  assign _zz_5018 = ($signed(data_mid_81_real) + $signed(_zz_421));
  assign _zz_5019 = _zz_5020;
  assign _zz_5020 = ($signed(_zz_5021) >>> _zz_424);
  assign _zz_5021 = _zz_5022;
  assign _zz_5022 = ($signed(data_mid_81_imag) + $signed(_zz_422));
  assign _zz_5023 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_86_real));
  assign _zz_5024 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_86_imag));
  assign _zz_5025 = fixTo_212_dout;
  assign _zz_5026 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_86_imag));
  assign _zz_5027 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_86_real));
  assign _zz_5028 = fixTo_213_dout;
  assign _zz_5029 = _zz_5030;
  assign _zz_5030 = ($signed(_zz_5031) >>> _zz_427);
  assign _zz_5031 = _zz_5032;
  assign _zz_5032 = ($signed(data_mid_84_real) - $signed(_zz_425));
  assign _zz_5033 = _zz_5034;
  assign _zz_5034 = ($signed(_zz_5035) >>> _zz_427);
  assign _zz_5035 = _zz_5036;
  assign _zz_5036 = ($signed(data_mid_84_imag) - $signed(_zz_426));
  assign _zz_5037 = _zz_5038;
  assign _zz_5038 = ($signed(_zz_5039) >>> _zz_428);
  assign _zz_5039 = _zz_5040;
  assign _zz_5040 = ($signed(data_mid_84_real) + $signed(_zz_425));
  assign _zz_5041 = _zz_5042;
  assign _zz_5042 = ($signed(_zz_5043) >>> _zz_428);
  assign _zz_5043 = _zz_5044;
  assign _zz_5044 = ($signed(data_mid_84_imag) + $signed(_zz_426));
  assign _zz_5045 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_87_real));
  assign _zz_5046 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_87_imag));
  assign _zz_5047 = fixTo_214_dout;
  assign _zz_5048 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_87_imag));
  assign _zz_5049 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_87_real));
  assign _zz_5050 = fixTo_215_dout;
  assign _zz_5051 = _zz_5052;
  assign _zz_5052 = ($signed(_zz_5053) >>> _zz_431);
  assign _zz_5053 = _zz_5054;
  assign _zz_5054 = ($signed(data_mid_85_real) - $signed(_zz_429));
  assign _zz_5055 = _zz_5056;
  assign _zz_5056 = ($signed(_zz_5057) >>> _zz_431);
  assign _zz_5057 = _zz_5058;
  assign _zz_5058 = ($signed(data_mid_85_imag) - $signed(_zz_430));
  assign _zz_5059 = _zz_5060;
  assign _zz_5060 = ($signed(_zz_5061) >>> _zz_432);
  assign _zz_5061 = _zz_5062;
  assign _zz_5062 = ($signed(data_mid_85_real) + $signed(_zz_429));
  assign _zz_5063 = _zz_5064;
  assign _zz_5064 = ($signed(_zz_5065) >>> _zz_432);
  assign _zz_5065 = _zz_5066;
  assign _zz_5066 = ($signed(data_mid_85_imag) + $signed(_zz_430));
  assign _zz_5067 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_90_real));
  assign _zz_5068 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_90_imag));
  assign _zz_5069 = fixTo_216_dout;
  assign _zz_5070 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_90_imag));
  assign _zz_5071 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_90_real));
  assign _zz_5072 = fixTo_217_dout;
  assign _zz_5073 = _zz_5074;
  assign _zz_5074 = ($signed(_zz_5075) >>> _zz_435);
  assign _zz_5075 = _zz_5076;
  assign _zz_5076 = ($signed(data_mid_88_real) - $signed(_zz_433));
  assign _zz_5077 = _zz_5078;
  assign _zz_5078 = ($signed(_zz_5079) >>> _zz_435);
  assign _zz_5079 = _zz_5080;
  assign _zz_5080 = ($signed(data_mid_88_imag) - $signed(_zz_434));
  assign _zz_5081 = _zz_5082;
  assign _zz_5082 = ($signed(_zz_5083) >>> _zz_436);
  assign _zz_5083 = _zz_5084;
  assign _zz_5084 = ($signed(data_mid_88_real) + $signed(_zz_433));
  assign _zz_5085 = _zz_5086;
  assign _zz_5086 = ($signed(_zz_5087) >>> _zz_436);
  assign _zz_5087 = _zz_5088;
  assign _zz_5088 = ($signed(data_mid_88_imag) + $signed(_zz_434));
  assign _zz_5089 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_91_real));
  assign _zz_5090 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_91_imag));
  assign _zz_5091 = fixTo_218_dout;
  assign _zz_5092 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_91_imag));
  assign _zz_5093 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_91_real));
  assign _zz_5094 = fixTo_219_dout;
  assign _zz_5095 = _zz_5096;
  assign _zz_5096 = ($signed(_zz_5097) >>> _zz_439);
  assign _zz_5097 = _zz_5098;
  assign _zz_5098 = ($signed(data_mid_89_real) - $signed(_zz_437));
  assign _zz_5099 = _zz_5100;
  assign _zz_5100 = ($signed(_zz_5101) >>> _zz_439);
  assign _zz_5101 = _zz_5102;
  assign _zz_5102 = ($signed(data_mid_89_imag) - $signed(_zz_438));
  assign _zz_5103 = _zz_5104;
  assign _zz_5104 = ($signed(_zz_5105) >>> _zz_440);
  assign _zz_5105 = _zz_5106;
  assign _zz_5106 = ($signed(data_mid_89_real) + $signed(_zz_437));
  assign _zz_5107 = _zz_5108;
  assign _zz_5108 = ($signed(_zz_5109) >>> _zz_440);
  assign _zz_5109 = _zz_5110;
  assign _zz_5110 = ($signed(data_mid_89_imag) + $signed(_zz_438));
  assign _zz_5111 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_94_real));
  assign _zz_5112 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_94_imag));
  assign _zz_5113 = fixTo_220_dout;
  assign _zz_5114 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_94_imag));
  assign _zz_5115 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_94_real));
  assign _zz_5116 = fixTo_221_dout;
  assign _zz_5117 = _zz_5118;
  assign _zz_5118 = ($signed(_zz_5119) >>> _zz_443);
  assign _zz_5119 = _zz_5120;
  assign _zz_5120 = ($signed(data_mid_92_real) - $signed(_zz_441));
  assign _zz_5121 = _zz_5122;
  assign _zz_5122 = ($signed(_zz_5123) >>> _zz_443);
  assign _zz_5123 = _zz_5124;
  assign _zz_5124 = ($signed(data_mid_92_imag) - $signed(_zz_442));
  assign _zz_5125 = _zz_5126;
  assign _zz_5126 = ($signed(_zz_5127) >>> _zz_444);
  assign _zz_5127 = _zz_5128;
  assign _zz_5128 = ($signed(data_mid_92_real) + $signed(_zz_441));
  assign _zz_5129 = _zz_5130;
  assign _zz_5130 = ($signed(_zz_5131) >>> _zz_444);
  assign _zz_5131 = _zz_5132;
  assign _zz_5132 = ($signed(data_mid_92_imag) + $signed(_zz_442));
  assign _zz_5133 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_95_real));
  assign _zz_5134 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_95_imag));
  assign _zz_5135 = fixTo_222_dout;
  assign _zz_5136 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_95_imag));
  assign _zz_5137 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_95_real));
  assign _zz_5138 = fixTo_223_dout;
  assign _zz_5139 = _zz_5140;
  assign _zz_5140 = ($signed(_zz_5141) >>> _zz_447);
  assign _zz_5141 = _zz_5142;
  assign _zz_5142 = ($signed(data_mid_93_real) - $signed(_zz_445));
  assign _zz_5143 = _zz_5144;
  assign _zz_5144 = ($signed(_zz_5145) >>> _zz_447);
  assign _zz_5145 = _zz_5146;
  assign _zz_5146 = ($signed(data_mid_93_imag) - $signed(_zz_446));
  assign _zz_5147 = _zz_5148;
  assign _zz_5148 = ($signed(_zz_5149) >>> _zz_448);
  assign _zz_5149 = _zz_5150;
  assign _zz_5150 = ($signed(data_mid_93_real) + $signed(_zz_445));
  assign _zz_5151 = _zz_5152;
  assign _zz_5152 = ($signed(_zz_5153) >>> _zz_448);
  assign _zz_5153 = _zz_5154;
  assign _zz_5154 = ($signed(data_mid_93_imag) + $signed(_zz_446));
  assign _zz_5155 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_98_real));
  assign _zz_5156 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_98_imag));
  assign _zz_5157 = fixTo_224_dout;
  assign _zz_5158 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_98_imag));
  assign _zz_5159 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_98_real));
  assign _zz_5160 = fixTo_225_dout;
  assign _zz_5161 = _zz_5162;
  assign _zz_5162 = ($signed(_zz_5163) >>> _zz_451);
  assign _zz_5163 = _zz_5164;
  assign _zz_5164 = ($signed(data_mid_96_real) - $signed(_zz_449));
  assign _zz_5165 = _zz_5166;
  assign _zz_5166 = ($signed(_zz_5167) >>> _zz_451);
  assign _zz_5167 = _zz_5168;
  assign _zz_5168 = ($signed(data_mid_96_imag) - $signed(_zz_450));
  assign _zz_5169 = _zz_5170;
  assign _zz_5170 = ($signed(_zz_5171) >>> _zz_452);
  assign _zz_5171 = _zz_5172;
  assign _zz_5172 = ($signed(data_mid_96_real) + $signed(_zz_449));
  assign _zz_5173 = _zz_5174;
  assign _zz_5174 = ($signed(_zz_5175) >>> _zz_452);
  assign _zz_5175 = _zz_5176;
  assign _zz_5176 = ($signed(data_mid_96_imag) + $signed(_zz_450));
  assign _zz_5177 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_99_real));
  assign _zz_5178 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_99_imag));
  assign _zz_5179 = fixTo_226_dout;
  assign _zz_5180 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_99_imag));
  assign _zz_5181 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_99_real));
  assign _zz_5182 = fixTo_227_dout;
  assign _zz_5183 = _zz_5184;
  assign _zz_5184 = ($signed(_zz_5185) >>> _zz_455);
  assign _zz_5185 = _zz_5186;
  assign _zz_5186 = ($signed(data_mid_97_real) - $signed(_zz_453));
  assign _zz_5187 = _zz_5188;
  assign _zz_5188 = ($signed(_zz_5189) >>> _zz_455);
  assign _zz_5189 = _zz_5190;
  assign _zz_5190 = ($signed(data_mid_97_imag) - $signed(_zz_454));
  assign _zz_5191 = _zz_5192;
  assign _zz_5192 = ($signed(_zz_5193) >>> _zz_456);
  assign _zz_5193 = _zz_5194;
  assign _zz_5194 = ($signed(data_mid_97_real) + $signed(_zz_453));
  assign _zz_5195 = _zz_5196;
  assign _zz_5196 = ($signed(_zz_5197) >>> _zz_456);
  assign _zz_5197 = _zz_5198;
  assign _zz_5198 = ($signed(data_mid_97_imag) + $signed(_zz_454));
  assign _zz_5199 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_102_real));
  assign _zz_5200 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_102_imag));
  assign _zz_5201 = fixTo_228_dout;
  assign _zz_5202 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_102_imag));
  assign _zz_5203 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_102_real));
  assign _zz_5204 = fixTo_229_dout;
  assign _zz_5205 = _zz_5206;
  assign _zz_5206 = ($signed(_zz_5207) >>> _zz_459);
  assign _zz_5207 = _zz_5208;
  assign _zz_5208 = ($signed(data_mid_100_real) - $signed(_zz_457));
  assign _zz_5209 = _zz_5210;
  assign _zz_5210 = ($signed(_zz_5211) >>> _zz_459);
  assign _zz_5211 = _zz_5212;
  assign _zz_5212 = ($signed(data_mid_100_imag) - $signed(_zz_458));
  assign _zz_5213 = _zz_5214;
  assign _zz_5214 = ($signed(_zz_5215) >>> _zz_460);
  assign _zz_5215 = _zz_5216;
  assign _zz_5216 = ($signed(data_mid_100_real) + $signed(_zz_457));
  assign _zz_5217 = _zz_5218;
  assign _zz_5218 = ($signed(_zz_5219) >>> _zz_460);
  assign _zz_5219 = _zz_5220;
  assign _zz_5220 = ($signed(data_mid_100_imag) + $signed(_zz_458));
  assign _zz_5221 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_103_real));
  assign _zz_5222 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_103_imag));
  assign _zz_5223 = fixTo_230_dout;
  assign _zz_5224 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_103_imag));
  assign _zz_5225 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_103_real));
  assign _zz_5226 = fixTo_231_dout;
  assign _zz_5227 = _zz_5228;
  assign _zz_5228 = ($signed(_zz_5229) >>> _zz_463);
  assign _zz_5229 = _zz_5230;
  assign _zz_5230 = ($signed(data_mid_101_real) - $signed(_zz_461));
  assign _zz_5231 = _zz_5232;
  assign _zz_5232 = ($signed(_zz_5233) >>> _zz_463);
  assign _zz_5233 = _zz_5234;
  assign _zz_5234 = ($signed(data_mid_101_imag) - $signed(_zz_462));
  assign _zz_5235 = _zz_5236;
  assign _zz_5236 = ($signed(_zz_5237) >>> _zz_464);
  assign _zz_5237 = _zz_5238;
  assign _zz_5238 = ($signed(data_mid_101_real) + $signed(_zz_461));
  assign _zz_5239 = _zz_5240;
  assign _zz_5240 = ($signed(_zz_5241) >>> _zz_464);
  assign _zz_5241 = _zz_5242;
  assign _zz_5242 = ($signed(data_mid_101_imag) + $signed(_zz_462));
  assign _zz_5243 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_106_real));
  assign _zz_5244 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_106_imag));
  assign _zz_5245 = fixTo_232_dout;
  assign _zz_5246 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_106_imag));
  assign _zz_5247 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_106_real));
  assign _zz_5248 = fixTo_233_dout;
  assign _zz_5249 = _zz_5250;
  assign _zz_5250 = ($signed(_zz_5251) >>> _zz_467);
  assign _zz_5251 = _zz_5252;
  assign _zz_5252 = ($signed(data_mid_104_real) - $signed(_zz_465));
  assign _zz_5253 = _zz_5254;
  assign _zz_5254 = ($signed(_zz_5255) >>> _zz_467);
  assign _zz_5255 = _zz_5256;
  assign _zz_5256 = ($signed(data_mid_104_imag) - $signed(_zz_466));
  assign _zz_5257 = _zz_5258;
  assign _zz_5258 = ($signed(_zz_5259) >>> _zz_468);
  assign _zz_5259 = _zz_5260;
  assign _zz_5260 = ($signed(data_mid_104_real) + $signed(_zz_465));
  assign _zz_5261 = _zz_5262;
  assign _zz_5262 = ($signed(_zz_5263) >>> _zz_468);
  assign _zz_5263 = _zz_5264;
  assign _zz_5264 = ($signed(data_mid_104_imag) + $signed(_zz_466));
  assign _zz_5265 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_107_real));
  assign _zz_5266 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_107_imag));
  assign _zz_5267 = fixTo_234_dout;
  assign _zz_5268 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_107_imag));
  assign _zz_5269 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_107_real));
  assign _zz_5270 = fixTo_235_dout;
  assign _zz_5271 = _zz_5272;
  assign _zz_5272 = ($signed(_zz_5273) >>> _zz_471);
  assign _zz_5273 = _zz_5274;
  assign _zz_5274 = ($signed(data_mid_105_real) - $signed(_zz_469));
  assign _zz_5275 = _zz_5276;
  assign _zz_5276 = ($signed(_zz_5277) >>> _zz_471);
  assign _zz_5277 = _zz_5278;
  assign _zz_5278 = ($signed(data_mid_105_imag) - $signed(_zz_470));
  assign _zz_5279 = _zz_5280;
  assign _zz_5280 = ($signed(_zz_5281) >>> _zz_472);
  assign _zz_5281 = _zz_5282;
  assign _zz_5282 = ($signed(data_mid_105_real) + $signed(_zz_469));
  assign _zz_5283 = _zz_5284;
  assign _zz_5284 = ($signed(_zz_5285) >>> _zz_472);
  assign _zz_5285 = _zz_5286;
  assign _zz_5286 = ($signed(data_mid_105_imag) + $signed(_zz_470));
  assign _zz_5287 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_110_real));
  assign _zz_5288 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_110_imag));
  assign _zz_5289 = fixTo_236_dout;
  assign _zz_5290 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_110_imag));
  assign _zz_5291 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_110_real));
  assign _zz_5292 = fixTo_237_dout;
  assign _zz_5293 = _zz_5294;
  assign _zz_5294 = ($signed(_zz_5295) >>> _zz_475);
  assign _zz_5295 = _zz_5296;
  assign _zz_5296 = ($signed(data_mid_108_real) - $signed(_zz_473));
  assign _zz_5297 = _zz_5298;
  assign _zz_5298 = ($signed(_zz_5299) >>> _zz_475);
  assign _zz_5299 = _zz_5300;
  assign _zz_5300 = ($signed(data_mid_108_imag) - $signed(_zz_474));
  assign _zz_5301 = _zz_5302;
  assign _zz_5302 = ($signed(_zz_5303) >>> _zz_476);
  assign _zz_5303 = _zz_5304;
  assign _zz_5304 = ($signed(data_mid_108_real) + $signed(_zz_473));
  assign _zz_5305 = _zz_5306;
  assign _zz_5306 = ($signed(_zz_5307) >>> _zz_476);
  assign _zz_5307 = _zz_5308;
  assign _zz_5308 = ($signed(data_mid_108_imag) + $signed(_zz_474));
  assign _zz_5309 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_111_real));
  assign _zz_5310 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_111_imag));
  assign _zz_5311 = fixTo_238_dout;
  assign _zz_5312 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_111_imag));
  assign _zz_5313 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_111_real));
  assign _zz_5314 = fixTo_239_dout;
  assign _zz_5315 = _zz_5316;
  assign _zz_5316 = ($signed(_zz_5317) >>> _zz_479);
  assign _zz_5317 = _zz_5318;
  assign _zz_5318 = ($signed(data_mid_109_real) - $signed(_zz_477));
  assign _zz_5319 = _zz_5320;
  assign _zz_5320 = ($signed(_zz_5321) >>> _zz_479);
  assign _zz_5321 = _zz_5322;
  assign _zz_5322 = ($signed(data_mid_109_imag) - $signed(_zz_478));
  assign _zz_5323 = _zz_5324;
  assign _zz_5324 = ($signed(_zz_5325) >>> _zz_480);
  assign _zz_5325 = _zz_5326;
  assign _zz_5326 = ($signed(data_mid_109_real) + $signed(_zz_477));
  assign _zz_5327 = _zz_5328;
  assign _zz_5328 = ($signed(_zz_5329) >>> _zz_480);
  assign _zz_5329 = _zz_5330;
  assign _zz_5330 = ($signed(data_mid_109_imag) + $signed(_zz_478));
  assign _zz_5331 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_114_real));
  assign _zz_5332 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_114_imag));
  assign _zz_5333 = fixTo_240_dout;
  assign _zz_5334 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_114_imag));
  assign _zz_5335 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_114_real));
  assign _zz_5336 = fixTo_241_dout;
  assign _zz_5337 = _zz_5338;
  assign _zz_5338 = ($signed(_zz_5339) >>> _zz_483);
  assign _zz_5339 = _zz_5340;
  assign _zz_5340 = ($signed(data_mid_112_real) - $signed(_zz_481));
  assign _zz_5341 = _zz_5342;
  assign _zz_5342 = ($signed(_zz_5343) >>> _zz_483);
  assign _zz_5343 = _zz_5344;
  assign _zz_5344 = ($signed(data_mid_112_imag) - $signed(_zz_482));
  assign _zz_5345 = _zz_5346;
  assign _zz_5346 = ($signed(_zz_5347) >>> _zz_484);
  assign _zz_5347 = _zz_5348;
  assign _zz_5348 = ($signed(data_mid_112_real) + $signed(_zz_481));
  assign _zz_5349 = _zz_5350;
  assign _zz_5350 = ($signed(_zz_5351) >>> _zz_484);
  assign _zz_5351 = _zz_5352;
  assign _zz_5352 = ($signed(data_mid_112_imag) + $signed(_zz_482));
  assign _zz_5353 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_115_real));
  assign _zz_5354 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_115_imag));
  assign _zz_5355 = fixTo_242_dout;
  assign _zz_5356 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_115_imag));
  assign _zz_5357 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_115_real));
  assign _zz_5358 = fixTo_243_dout;
  assign _zz_5359 = _zz_5360;
  assign _zz_5360 = ($signed(_zz_5361) >>> _zz_487);
  assign _zz_5361 = _zz_5362;
  assign _zz_5362 = ($signed(data_mid_113_real) - $signed(_zz_485));
  assign _zz_5363 = _zz_5364;
  assign _zz_5364 = ($signed(_zz_5365) >>> _zz_487);
  assign _zz_5365 = _zz_5366;
  assign _zz_5366 = ($signed(data_mid_113_imag) - $signed(_zz_486));
  assign _zz_5367 = _zz_5368;
  assign _zz_5368 = ($signed(_zz_5369) >>> _zz_488);
  assign _zz_5369 = _zz_5370;
  assign _zz_5370 = ($signed(data_mid_113_real) + $signed(_zz_485));
  assign _zz_5371 = _zz_5372;
  assign _zz_5372 = ($signed(_zz_5373) >>> _zz_488);
  assign _zz_5373 = _zz_5374;
  assign _zz_5374 = ($signed(data_mid_113_imag) + $signed(_zz_486));
  assign _zz_5375 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_118_real));
  assign _zz_5376 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_118_imag));
  assign _zz_5377 = fixTo_244_dout;
  assign _zz_5378 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_118_imag));
  assign _zz_5379 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_118_real));
  assign _zz_5380 = fixTo_245_dout;
  assign _zz_5381 = _zz_5382;
  assign _zz_5382 = ($signed(_zz_5383) >>> _zz_491);
  assign _zz_5383 = _zz_5384;
  assign _zz_5384 = ($signed(data_mid_116_real) - $signed(_zz_489));
  assign _zz_5385 = _zz_5386;
  assign _zz_5386 = ($signed(_zz_5387) >>> _zz_491);
  assign _zz_5387 = _zz_5388;
  assign _zz_5388 = ($signed(data_mid_116_imag) - $signed(_zz_490));
  assign _zz_5389 = _zz_5390;
  assign _zz_5390 = ($signed(_zz_5391) >>> _zz_492);
  assign _zz_5391 = _zz_5392;
  assign _zz_5392 = ($signed(data_mid_116_real) + $signed(_zz_489));
  assign _zz_5393 = _zz_5394;
  assign _zz_5394 = ($signed(_zz_5395) >>> _zz_492);
  assign _zz_5395 = _zz_5396;
  assign _zz_5396 = ($signed(data_mid_116_imag) + $signed(_zz_490));
  assign _zz_5397 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_119_real));
  assign _zz_5398 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_119_imag));
  assign _zz_5399 = fixTo_246_dout;
  assign _zz_5400 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_119_imag));
  assign _zz_5401 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_119_real));
  assign _zz_5402 = fixTo_247_dout;
  assign _zz_5403 = _zz_5404;
  assign _zz_5404 = ($signed(_zz_5405) >>> _zz_495);
  assign _zz_5405 = _zz_5406;
  assign _zz_5406 = ($signed(data_mid_117_real) - $signed(_zz_493));
  assign _zz_5407 = _zz_5408;
  assign _zz_5408 = ($signed(_zz_5409) >>> _zz_495);
  assign _zz_5409 = _zz_5410;
  assign _zz_5410 = ($signed(data_mid_117_imag) - $signed(_zz_494));
  assign _zz_5411 = _zz_5412;
  assign _zz_5412 = ($signed(_zz_5413) >>> _zz_496);
  assign _zz_5413 = _zz_5414;
  assign _zz_5414 = ($signed(data_mid_117_real) + $signed(_zz_493));
  assign _zz_5415 = _zz_5416;
  assign _zz_5416 = ($signed(_zz_5417) >>> _zz_496);
  assign _zz_5417 = _zz_5418;
  assign _zz_5418 = ($signed(data_mid_117_imag) + $signed(_zz_494));
  assign _zz_5419 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_122_real));
  assign _zz_5420 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_122_imag));
  assign _zz_5421 = fixTo_248_dout;
  assign _zz_5422 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_122_imag));
  assign _zz_5423 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_122_real));
  assign _zz_5424 = fixTo_249_dout;
  assign _zz_5425 = _zz_5426;
  assign _zz_5426 = ($signed(_zz_5427) >>> _zz_499);
  assign _zz_5427 = _zz_5428;
  assign _zz_5428 = ($signed(data_mid_120_real) - $signed(_zz_497));
  assign _zz_5429 = _zz_5430;
  assign _zz_5430 = ($signed(_zz_5431) >>> _zz_499);
  assign _zz_5431 = _zz_5432;
  assign _zz_5432 = ($signed(data_mid_120_imag) - $signed(_zz_498));
  assign _zz_5433 = _zz_5434;
  assign _zz_5434 = ($signed(_zz_5435) >>> _zz_500);
  assign _zz_5435 = _zz_5436;
  assign _zz_5436 = ($signed(data_mid_120_real) + $signed(_zz_497));
  assign _zz_5437 = _zz_5438;
  assign _zz_5438 = ($signed(_zz_5439) >>> _zz_500);
  assign _zz_5439 = _zz_5440;
  assign _zz_5440 = ($signed(data_mid_120_imag) + $signed(_zz_498));
  assign _zz_5441 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_123_real));
  assign _zz_5442 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_123_imag));
  assign _zz_5443 = fixTo_250_dout;
  assign _zz_5444 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_123_imag));
  assign _zz_5445 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_123_real));
  assign _zz_5446 = fixTo_251_dout;
  assign _zz_5447 = _zz_5448;
  assign _zz_5448 = ($signed(_zz_5449) >>> _zz_503);
  assign _zz_5449 = _zz_5450;
  assign _zz_5450 = ($signed(data_mid_121_real) - $signed(_zz_501));
  assign _zz_5451 = _zz_5452;
  assign _zz_5452 = ($signed(_zz_5453) >>> _zz_503);
  assign _zz_5453 = _zz_5454;
  assign _zz_5454 = ($signed(data_mid_121_imag) - $signed(_zz_502));
  assign _zz_5455 = _zz_5456;
  assign _zz_5456 = ($signed(_zz_5457) >>> _zz_504);
  assign _zz_5457 = _zz_5458;
  assign _zz_5458 = ($signed(data_mid_121_real) + $signed(_zz_501));
  assign _zz_5459 = _zz_5460;
  assign _zz_5460 = ($signed(_zz_5461) >>> _zz_504);
  assign _zz_5461 = _zz_5462;
  assign _zz_5462 = ($signed(data_mid_121_imag) + $signed(_zz_502));
  assign _zz_5463 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_126_real));
  assign _zz_5464 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_126_imag));
  assign _zz_5465 = fixTo_252_dout;
  assign _zz_5466 = ($signed(twiddle_factor_table_1_real) * $signed(data_mid_126_imag));
  assign _zz_5467 = ($signed(twiddle_factor_table_1_imag) * $signed(data_mid_126_real));
  assign _zz_5468 = fixTo_253_dout;
  assign _zz_5469 = _zz_5470;
  assign _zz_5470 = ($signed(_zz_5471) >>> _zz_507);
  assign _zz_5471 = _zz_5472;
  assign _zz_5472 = ($signed(data_mid_124_real) - $signed(_zz_505));
  assign _zz_5473 = _zz_5474;
  assign _zz_5474 = ($signed(_zz_5475) >>> _zz_507);
  assign _zz_5475 = _zz_5476;
  assign _zz_5476 = ($signed(data_mid_124_imag) - $signed(_zz_506));
  assign _zz_5477 = _zz_5478;
  assign _zz_5478 = ($signed(_zz_5479) >>> _zz_508);
  assign _zz_5479 = _zz_5480;
  assign _zz_5480 = ($signed(data_mid_124_real) + $signed(_zz_505));
  assign _zz_5481 = _zz_5482;
  assign _zz_5482 = ($signed(_zz_5483) >>> _zz_508);
  assign _zz_5483 = _zz_5484;
  assign _zz_5484 = ($signed(data_mid_124_imag) + $signed(_zz_506));
  assign _zz_5485 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_127_real));
  assign _zz_5486 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_127_imag));
  assign _zz_5487 = fixTo_254_dout;
  assign _zz_5488 = ($signed(twiddle_factor_table_2_real) * $signed(data_mid_127_imag));
  assign _zz_5489 = ($signed(twiddle_factor_table_2_imag) * $signed(data_mid_127_real));
  assign _zz_5490 = fixTo_255_dout;
  assign _zz_5491 = _zz_5492;
  assign _zz_5492 = ($signed(_zz_5493) >>> _zz_511);
  assign _zz_5493 = _zz_5494;
  assign _zz_5494 = ($signed(data_mid_125_real) - $signed(_zz_509));
  assign _zz_5495 = _zz_5496;
  assign _zz_5496 = ($signed(_zz_5497) >>> _zz_511);
  assign _zz_5497 = _zz_5498;
  assign _zz_5498 = ($signed(data_mid_125_imag) - $signed(_zz_510));
  assign _zz_5499 = _zz_5500;
  assign _zz_5500 = ($signed(_zz_5501) >>> _zz_512);
  assign _zz_5501 = _zz_5502;
  assign _zz_5502 = ($signed(data_mid_125_real) + $signed(_zz_509));
  assign _zz_5503 = _zz_5504;
  assign _zz_5504 = ($signed(_zz_5505) >>> _zz_512);
  assign _zz_5505 = _zz_5506;
  assign _zz_5506 = ($signed(data_mid_125_imag) + $signed(_zz_510));
  assign _zz_5507 = ($signed(twiddle_factor_table_3_real) * $signed(data_mid_4_real));
  assign _zz_5508 = ($signed(twiddle_factor_table_3_imag) * $signed(data_mid_4_imag));
  assign _zz_5509 = fixTo_256_dout;
  assign _zz_5510 = ($signed(twiddle_factor_table_3_real) * $signed(data_mid_4_imag));
  assign _zz_5511 = ($signed(twiddle_factor_table_3_imag) * $signed(data_mid_4_real));
  assign _zz_5512 = fixTo_257_dout;
  assign _zz_5513 = _zz_5514;
  assign _zz_5514 = ($signed(_zz_5515) >>> _zz_515);
  assign _zz_5515 = _zz_5516;
  assign _zz_5516 = ($signed(data_mid_0_real) - $signed(_zz_513));
  assign _zz_5517 = _zz_5518;
  assign _zz_5518 = ($signed(_zz_5519) >>> _zz_515);
  assign _zz_5519 = _zz_5520;
  assign _zz_5520 = ($signed(data_mid_0_imag) - $signed(_zz_514));
  assign _zz_5521 = _zz_5522;
  assign _zz_5522 = ($signed(_zz_5523) >>> _zz_516);
  assign _zz_5523 = _zz_5524;
  assign _zz_5524 = ($signed(data_mid_0_real) + $signed(_zz_513));
  assign _zz_5525 = _zz_5526;
  assign _zz_5526 = ($signed(_zz_5527) >>> _zz_516);
  assign _zz_5527 = _zz_5528;
  assign _zz_5528 = ($signed(data_mid_0_imag) + $signed(_zz_514));
  assign _zz_5529 = ($signed(twiddle_factor_table_4_real) * $signed(data_mid_5_real));
  assign _zz_5530 = ($signed(twiddle_factor_table_4_imag) * $signed(data_mid_5_imag));
  assign _zz_5531 = fixTo_258_dout;
  assign _zz_5532 = ($signed(twiddle_factor_table_4_real) * $signed(data_mid_5_imag));
  assign _zz_5533 = ($signed(twiddle_factor_table_4_imag) * $signed(data_mid_5_real));
  assign _zz_5534 = fixTo_259_dout;
  assign _zz_5535 = _zz_5536;
  assign _zz_5536 = ($signed(_zz_5537) >>> _zz_519);
  assign _zz_5537 = _zz_5538;
  assign _zz_5538 = ($signed(data_mid_1_real) - $signed(_zz_517));
  assign _zz_5539 = _zz_5540;
  assign _zz_5540 = ($signed(_zz_5541) >>> _zz_519);
  assign _zz_5541 = _zz_5542;
  assign _zz_5542 = ($signed(data_mid_1_imag) - $signed(_zz_518));
  assign _zz_5543 = _zz_5544;
  assign _zz_5544 = ($signed(_zz_5545) >>> _zz_520);
  assign _zz_5545 = _zz_5546;
  assign _zz_5546 = ($signed(data_mid_1_real) + $signed(_zz_517));
  assign _zz_5547 = _zz_5548;
  assign _zz_5548 = ($signed(_zz_5549) >>> _zz_520);
  assign _zz_5549 = _zz_5550;
  assign _zz_5550 = ($signed(data_mid_1_imag) + $signed(_zz_518));
  assign _zz_5551 = ($signed(twiddle_factor_table_5_real) * $signed(data_mid_6_real));
  assign _zz_5552 = ($signed(twiddle_factor_table_5_imag) * $signed(data_mid_6_imag));
  assign _zz_5553 = fixTo_260_dout;
  assign _zz_5554 = ($signed(twiddle_factor_table_5_real) * $signed(data_mid_6_imag));
  assign _zz_5555 = ($signed(twiddle_factor_table_5_imag) * $signed(data_mid_6_real));
  assign _zz_5556 = fixTo_261_dout;
  assign _zz_5557 = _zz_5558;
  assign _zz_5558 = ($signed(_zz_5559) >>> _zz_523);
  assign _zz_5559 = _zz_5560;
  assign _zz_5560 = ($signed(data_mid_2_real) - $signed(_zz_521));
  assign _zz_5561 = _zz_5562;
  assign _zz_5562 = ($signed(_zz_5563) >>> _zz_523);
  assign _zz_5563 = _zz_5564;
  assign _zz_5564 = ($signed(data_mid_2_imag) - $signed(_zz_522));
  assign _zz_5565 = _zz_5566;
  assign _zz_5566 = ($signed(_zz_5567) >>> _zz_524);
  assign _zz_5567 = _zz_5568;
  assign _zz_5568 = ($signed(data_mid_2_real) + $signed(_zz_521));
  assign _zz_5569 = _zz_5570;
  assign _zz_5570 = ($signed(_zz_5571) >>> _zz_524);
  assign _zz_5571 = _zz_5572;
  assign _zz_5572 = ($signed(data_mid_2_imag) + $signed(_zz_522));
  assign _zz_5573 = ($signed(twiddle_factor_table_6_real) * $signed(data_mid_7_real));
  assign _zz_5574 = ($signed(twiddle_factor_table_6_imag) * $signed(data_mid_7_imag));
  assign _zz_5575 = fixTo_262_dout;
  assign _zz_5576 = ($signed(twiddle_factor_table_6_real) * $signed(data_mid_7_imag));
  assign _zz_5577 = ($signed(twiddle_factor_table_6_imag) * $signed(data_mid_7_real));
  assign _zz_5578 = fixTo_263_dout;
  assign _zz_5579 = _zz_5580;
  assign _zz_5580 = ($signed(_zz_5581) >>> _zz_527);
  assign _zz_5581 = _zz_5582;
  assign _zz_5582 = ($signed(data_mid_3_real) - $signed(_zz_525));
  assign _zz_5583 = _zz_5584;
  assign _zz_5584 = ($signed(_zz_5585) >>> _zz_527);
  assign _zz_5585 = _zz_5586;
  assign _zz_5586 = ($signed(data_mid_3_imag) - $signed(_zz_526));
  assign _zz_5587 = _zz_5588;
  assign _zz_5588 = ($signed(_zz_5589) >>> _zz_528);
  assign _zz_5589 = _zz_5590;
  assign _zz_5590 = ($signed(data_mid_3_real) + $signed(_zz_525));
  assign _zz_5591 = _zz_5592;
  assign _zz_5592 = ($signed(_zz_5593) >>> _zz_528);
  assign _zz_5593 = _zz_5594;
  assign _zz_5594 = ($signed(data_mid_3_imag) + $signed(_zz_526));
  assign _zz_5595 = ($signed(twiddle_factor_table_3_real) * $signed(data_mid_12_real));
  assign _zz_5596 = ($signed(twiddle_factor_table_3_imag) * $signed(data_mid_12_imag));
  assign _zz_5597 = fixTo_264_dout;
  assign _zz_5598 = ($signed(twiddle_factor_table_3_real) * $signed(data_mid_12_imag));
  assign _zz_5599 = ($signed(twiddle_factor_table_3_imag) * $signed(data_mid_12_real));
  assign _zz_5600 = fixTo_265_dout;
  assign _zz_5601 = _zz_5602;
  assign _zz_5602 = ($signed(_zz_5603) >>> _zz_531);
  assign _zz_5603 = _zz_5604;
  assign _zz_5604 = ($signed(data_mid_8_real) - $signed(_zz_529));
  assign _zz_5605 = _zz_5606;
  assign _zz_5606 = ($signed(_zz_5607) >>> _zz_531);
  assign _zz_5607 = _zz_5608;
  assign _zz_5608 = ($signed(data_mid_8_imag) - $signed(_zz_530));
  assign _zz_5609 = _zz_5610;
  assign _zz_5610 = ($signed(_zz_5611) >>> _zz_532);
  assign _zz_5611 = _zz_5612;
  assign _zz_5612 = ($signed(data_mid_8_real) + $signed(_zz_529));
  assign _zz_5613 = _zz_5614;
  assign _zz_5614 = ($signed(_zz_5615) >>> _zz_532);
  assign _zz_5615 = _zz_5616;
  assign _zz_5616 = ($signed(data_mid_8_imag) + $signed(_zz_530));
  assign _zz_5617 = ($signed(twiddle_factor_table_4_real) * $signed(data_mid_13_real));
  assign _zz_5618 = ($signed(twiddle_factor_table_4_imag) * $signed(data_mid_13_imag));
  assign _zz_5619 = fixTo_266_dout;
  assign _zz_5620 = ($signed(twiddle_factor_table_4_real) * $signed(data_mid_13_imag));
  assign _zz_5621 = ($signed(twiddle_factor_table_4_imag) * $signed(data_mid_13_real));
  assign _zz_5622 = fixTo_267_dout;
  assign _zz_5623 = _zz_5624;
  assign _zz_5624 = ($signed(_zz_5625) >>> _zz_535);
  assign _zz_5625 = _zz_5626;
  assign _zz_5626 = ($signed(data_mid_9_real) - $signed(_zz_533));
  assign _zz_5627 = _zz_5628;
  assign _zz_5628 = ($signed(_zz_5629) >>> _zz_535);
  assign _zz_5629 = _zz_5630;
  assign _zz_5630 = ($signed(data_mid_9_imag) - $signed(_zz_534));
  assign _zz_5631 = _zz_5632;
  assign _zz_5632 = ($signed(_zz_5633) >>> _zz_536);
  assign _zz_5633 = _zz_5634;
  assign _zz_5634 = ($signed(data_mid_9_real) + $signed(_zz_533));
  assign _zz_5635 = _zz_5636;
  assign _zz_5636 = ($signed(_zz_5637) >>> _zz_536);
  assign _zz_5637 = _zz_5638;
  assign _zz_5638 = ($signed(data_mid_9_imag) + $signed(_zz_534));
  assign _zz_5639 = ($signed(twiddle_factor_table_5_real) * $signed(data_mid_14_real));
  assign _zz_5640 = ($signed(twiddle_factor_table_5_imag) * $signed(data_mid_14_imag));
  assign _zz_5641 = fixTo_268_dout;
  assign _zz_5642 = ($signed(twiddle_factor_table_5_real) * $signed(data_mid_14_imag));
  assign _zz_5643 = ($signed(twiddle_factor_table_5_imag) * $signed(data_mid_14_real));
  assign _zz_5644 = fixTo_269_dout;
  assign _zz_5645 = _zz_5646;
  assign _zz_5646 = ($signed(_zz_5647) >>> _zz_539);
  assign _zz_5647 = _zz_5648;
  assign _zz_5648 = ($signed(data_mid_10_real) - $signed(_zz_537));
  assign _zz_5649 = _zz_5650;
  assign _zz_5650 = ($signed(_zz_5651) >>> _zz_539);
  assign _zz_5651 = _zz_5652;
  assign _zz_5652 = ($signed(data_mid_10_imag) - $signed(_zz_538));
  assign _zz_5653 = _zz_5654;
  assign _zz_5654 = ($signed(_zz_5655) >>> _zz_540);
  assign _zz_5655 = _zz_5656;
  assign _zz_5656 = ($signed(data_mid_10_real) + $signed(_zz_537));
  assign _zz_5657 = _zz_5658;
  assign _zz_5658 = ($signed(_zz_5659) >>> _zz_540);
  assign _zz_5659 = _zz_5660;
  assign _zz_5660 = ($signed(data_mid_10_imag) + $signed(_zz_538));
  assign _zz_5661 = ($signed(twiddle_factor_table_6_real) * $signed(data_mid_15_real));
  assign _zz_5662 = ($signed(twiddle_factor_table_6_imag) * $signed(data_mid_15_imag));
  assign _zz_5663 = fixTo_270_dout;
  assign _zz_5664 = ($signed(twiddle_factor_table_6_real) * $signed(data_mid_15_imag));
  assign _zz_5665 = ($signed(twiddle_factor_table_6_imag) * $signed(data_mid_15_real));
  assign _zz_5666 = fixTo_271_dout;
  assign _zz_5667 = _zz_5668;
  assign _zz_5668 = ($signed(_zz_5669) >>> _zz_543);
  assign _zz_5669 = _zz_5670;
  assign _zz_5670 = ($signed(data_mid_11_real) - $signed(_zz_541));
  assign _zz_5671 = _zz_5672;
  assign _zz_5672 = ($signed(_zz_5673) >>> _zz_543);
  assign _zz_5673 = _zz_5674;
  assign _zz_5674 = ($signed(data_mid_11_imag) - $signed(_zz_542));
  assign _zz_5675 = _zz_5676;
  assign _zz_5676 = ($signed(_zz_5677) >>> _zz_544);
  assign _zz_5677 = _zz_5678;
  assign _zz_5678 = ($signed(data_mid_11_real) + $signed(_zz_541));
  assign _zz_5679 = _zz_5680;
  assign _zz_5680 = ($signed(_zz_5681) >>> _zz_544);
  assign _zz_5681 = _zz_5682;
  assign _zz_5682 = ($signed(data_mid_11_imag) + $signed(_zz_542));
  assign _zz_5683 = ($signed(twiddle_factor_table_3_real) * $signed(data_mid_20_real));
  assign _zz_5684 = ($signed(twiddle_factor_table_3_imag) * $signed(data_mid_20_imag));
  assign _zz_5685 = fixTo_272_dout;
  assign _zz_5686 = ($signed(twiddle_factor_table_3_real) * $signed(data_mid_20_imag));
  assign _zz_5687 = ($signed(twiddle_factor_table_3_imag) * $signed(data_mid_20_real));
  assign _zz_5688 = fixTo_273_dout;
  assign _zz_5689 = _zz_5690;
  assign _zz_5690 = ($signed(_zz_5691) >>> _zz_547);
  assign _zz_5691 = _zz_5692;
  assign _zz_5692 = ($signed(data_mid_16_real) - $signed(_zz_545));
  assign _zz_5693 = _zz_5694;
  assign _zz_5694 = ($signed(_zz_5695) >>> _zz_547);
  assign _zz_5695 = _zz_5696;
  assign _zz_5696 = ($signed(data_mid_16_imag) - $signed(_zz_546));
  assign _zz_5697 = _zz_5698;
  assign _zz_5698 = ($signed(_zz_5699) >>> _zz_548);
  assign _zz_5699 = _zz_5700;
  assign _zz_5700 = ($signed(data_mid_16_real) + $signed(_zz_545));
  assign _zz_5701 = _zz_5702;
  assign _zz_5702 = ($signed(_zz_5703) >>> _zz_548);
  assign _zz_5703 = _zz_5704;
  assign _zz_5704 = ($signed(data_mid_16_imag) + $signed(_zz_546));
  assign _zz_5705 = ($signed(twiddle_factor_table_4_real) * $signed(data_mid_21_real));
  assign _zz_5706 = ($signed(twiddle_factor_table_4_imag) * $signed(data_mid_21_imag));
  assign _zz_5707 = fixTo_274_dout;
  assign _zz_5708 = ($signed(twiddle_factor_table_4_real) * $signed(data_mid_21_imag));
  assign _zz_5709 = ($signed(twiddle_factor_table_4_imag) * $signed(data_mid_21_real));
  assign _zz_5710 = fixTo_275_dout;
  assign _zz_5711 = _zz_5712;
  assign _zz_5712 = ($signed(_zz_5713) >>> _zz_551);
  assign _zz_5713 = _zz_5714;
  assign _zz_5714 = ($signed(data_mid_17_real) - $signed(_zz_549));
  assign _zz_5715 = _zz_5716;
  assign _zz_5716 = ($signed(_zz_5717) >>> _zz_551);
  assign _zz_5717 = _zz_5718;
  assign _zz_5718 = ($signed(data_mid_17_imag) - $signed(_zz_550));
  assign _zz_5719 = _zz_5720;
  assign _zz_5720 = ($signed(_zz_5721) >>> _zz_552);
  assign _zz_5721 = _zz_5722;
  assign _zz_5722 = ($signed(data_mid_17_real) + $signed(_zz_549));
  assign _zz_5723 = _zz_5724;
  assign _zz_5724 = ($signed(_zz_5725) >>> _zz_552);
  assign _zz_5725 = _zz_5726;
  assign _zz_5726 = ($signed(data_mid_17_imag) + $signed(_zz_550));
  assign _zz_5727 = ($signed(twiddle_factor_table_5_real) * $signed(data_mid_22_real));
  assign _zz_5728 = ($signed(twiddle_factor_table_5_imag) * $signed(data_mid_22_imag));
  assign _zz_5729 = fixTo_276_dout;
  assign _zz_5730 = ($signed(twiddle_factor_table_5_real) * $signed(data_mid_22_imag));
  assign _zz_5731 = ($signed(twiddle_factor_table_5_imag) * $signed(data_mid_22_real));
  assign _zz_5732 = fixTo_277_dout;
  assign _zz_5733 = _zz_5734;
  assign _zz_5734 = ($signed(_zz_5735) >>> _zz_555);
  assign _zz_5735 = _zz_5736;
  assign _zz_5736 = ($signed(data_mid_18_real) - $signed(_zz_553));
  assign _zz_5737 = _zz_5738;
  assign _zz_5738 = ($signed(_zz_5739) >>> _zz_555);
  assign _zz_5739 = _zz_5740;
  assign _zz_5740 = ($signed(data_mid_18_imag) - $signed(_zz_554));
  assign _zz_5741 = _zz_5742;
  assign _zz_5742 = ($signed(_zz_5743) >>> _zz_556);
  assign _zz_5743 = _zz_5744;
  assign _zz_5744 = ($signed(data_mid_18_real) + $signed(_zz_553));
  assign _zz_5745 = _zz_5746;
  assign _zz_5746 = ($signed(_zz_5747) >>> _zz_556);
  assign _zz_5747 = _zz_5748;
  assign _zz_5748 = ($signed(data_mid_18_imag) + $signed(_zz_554));
  assign _zz_5749 = ($signed(twiddle_factor_table_6_real) * $signed(data_mid_23_real));
  assign _zz_5750 = ($signed(twiddle_factor_table_6_imag) * $signed(data_mid_23_imag));
  assign _zz_5751 = fixTo_278_dout;
  assign _zz_5752 = ($signed(twiddle_factor_table_6_real) * $signed(data_mid_23_imag));
  assign _zz_5753 = ($signed(twiddle_factor_table_6_imag) * $signed(data_mid_23_real));
  assign _zz_5754 = fixTo_279_dout;
  assign _zz_5755 = _zz_5756;
  assign _zz_5756 = ($signed(_zz_5757) >>> _zz_559);
  assign _zz_5757 = _zz_5758;
  assign _zz_5758 = ($signed(data_mid_19_real) - $signed(_zz_557));
  assign _zz_5759 = _zz_5760;
  assign _zz_5760 = ($signed(_zz_5761) >>> _zz_559);
  assign _zz_5761 = _zz_5762;
  assign _zz_5762 = ($signed(data_mid_19_imag) - $signed(_zz_558));
  assign _zz_5763 = _zz_5764;
  assign _zz_5764 = ($signed(_zz_5765) >>> _zz_560);
  assign _zz_5765 = _zz_5766;
  assign _zz_5766 = ($signed(data_mid_19_real) + $signed(_zz_557));
  assign _zz_5767 = _zz_5768;
  assign _zz_5768 = ($signed(_zz_5769) >>> _zz_560);
  assign _zz_5769 = _zz_5770;
  assign _zz_5770 = ($signed(data_mid_19_imag) + $signed(_zz_558));
  assign _zz_5771 = ($signed(twiddle_factor_table_3_real) * $signed(data_mid_28_real));
  assign _zz_5772 = ($signed(twiddle_factor_table_3_imag) * $signed(data_mid_28_imag));
  assign _zz_5773 = fixTo_280_dout;
  assign _zz_5774 = ($signed(twiddle_factor_table_3_real) * $signed(data_mid_28_imag));
  assign _zz_5775 = ($signed(twiddle_factor_table_3_imag) * $signed(data_mid_28_real));
  assign _zz_5776 = fixTo_281_dout;
  assign _zz_5777 = _zz_5778;
  assign _zz_5778 = ($signed(_zz_5779) >>> _zz_563);
  assign _zz_5779 = _zz_5780;
  assign _zz_5780 = ($signed(data_mid_24_real) - $signed(_zz_561));
  assign _zz_5781 = _zz_5782;
  assign _zz_5782 = ($signed(_zz_5783) >>> _zz_563);
  assign _zz_5783 = _zz_5784;
  assign _zz_5784 = ($signed(data_mid_24_imag) - $signed(_zz_562));
  assign _zz_5785 = _zz_5786;
  assign _zz_5786 = ($signed(_zz_5787) >>> _zz_564);
  assign _zz_5787 = _zz_5788;
  assign _zz_5788 = ($signed(data_mid_24_real) + $signed(_zz_561));
  assign _zz_5789 = _zz_5790;
  assign _zz_5790 = ($signed(_zz_5791) >>> _zz_564);
  assign _zz_5791 = _zz_5792;
  assign _zz_5792 = ($signed(data_mid_24_imag) + $signed(_zz_562));
  assign _zz_5793 = ($signed(twiddle_factor_table_4_real) * $signed(data_mid_29_real));
  assign _zz_5794 = ($signed(twiddle_factor_table_4_imag) * $signed(data_mid_29_imag));
  assign _zz_5795 = fixTo_282_dout;
  assign _zz_5796 = ($signed(twiddle_factor_table_4_real) * $signed(data_mid_29_imag));
  assign _zz_5797 = ($signed(twiddle_factor_table_4_imag) * $signed(data_mid_29_real));
  assign _zz_5798 = fixTo_283_dout;
  assign _zz_5799 = _zz_5800;
  assign _zz_5800 = ($signed(_zz_5801) >>> _zz_567);
  assign _zz_5801 = _zz_5802;
  assign _zz_5802 = ($signed(data_mid_25_real) - $signed(_zz_565));
  assign _zz_5803 = _zz_5804;
  assign _zz_5804 = ($signed(_zz_5805) >>> _zz_567);
  assign _zz_5805 = _zz_5806;
  assign _zz_5806 = ($signed(data_mid_25_imag) - $signed(_zz_566));
  assign _zz_5807 = _zz_5808;
  assign _zz_5808 = ($signed(_zz_5809) >>> _zz_568);
  assign _zz_5809 = _zz_5810;
  assign _zz_5810 = ($signed(data_mid_25_real) + $signed(_zz_565));
  assign _zz_5811 = _zz_5812;
  assign _zz_5812 = ($signed(_zz_5813) >>> _zz_568);
  assign _zz_5813 = _zz_5814;
  assign _zz_5814 = ($signed(data_mid_25_imag) + $signed(_zz_566));
  assign _zz_5815 = ($signed(twiddle_factor_table_5_real) * $signed(data_mid_30_real));
  assign _zz_5816 = ($signed(twiddle_factor_table_5_imag) * $signed(data_mid_30_imag));
  assign _zz_5817 = fixTo_284_dout;
  assign _zz_5818 = ($signed(twiddle_factor_table_5_real) * $signed(data_mid_30_imag));
  assign _zz_5819 = ($signed(twiddle_factor_table_5_imag) * $signed(data_mid_30_real));
  assign _zz_5820 = fixTo_285_dout;
  assign _zz_5821 = _zz_5822;
  assign _zz_5822 = ($signed(_zz_5823) >>> _zz_571);
  assign _zz_5823 = _zz_5824;
  assign _zz_5824 = ($signed(data_mid_26_real) - $signed(_zz_569));
  assign _zz_5825 = _zz_5826;
  assign _zz_5826 = ($signed(_zz_5827) >>> _zz_571);
  assign _zz_5827 = _zz_5828;
  assign _zz_5828 = ($signed(data_mid_26_imag) - $signed(_zz_570));
  assign _zz_5829 = _zz_5830;
  assign _zz_5830 = ($signed(_zz_5831) >>> _zz_572);
  assign _zz_5831 = _zz_5832;
  assign _zz_5832 = ($signed(data_mid_26_real) + $signed(_zz_569));
  assign _zz_5833 = _zz_5834;
  assign _zz_5834 = ($signed(_zz_5835) >>> _zz_572);
  assign _zz_5835 = _zz_5836;
  assign _zz_5836 = ($signed(data_mid_26_imag) + $signed(_zz_570));
  assign _zz_5837 = ($signed(twiddle_factor_table_6_real) * $signed(data_mid_31_real));
  assign _zz_5838 = ($signed(twiddle_factor_table_6_imag) * $signed(data_mid_31_imag));
  assign _zz_5839 = fixTo_286_dout;
  assign _zz_5840 = ($signed(twiddle_factor_table_6_real) * $signed(data_mid_31_imag));
  assign _zz_5841 = ($signed(twiddle_factor_table_6_imag) * $signed(data_mid_31_real));
  assign _zz_5842 = fixTo_287_dout;
  assign _zz_5843 = _zz_5844;
  assign _zz_5844 = ($signed(_zz_5845) >>> _zz_575);
  assign _zz_5845 = _zz_5846;
  assign _zz_5846 = ($signed(data_mid_27_real) - $signed(_zz_573));
  assign _zz_5847 = _zz_5848;
  assign _zz_5848 = ($signed(_zz_5849) >>> _zz_575);
  assign _zz_5849 = _zz_5850;
  assign _zz_5850 = ($signed(data_mid_27_imag) - $signed(_zz_574));
  assign _zz_5851 = _zz_5852;
  assign _zz_5852 = ($signed(_zz_5853) >>> _zz_576);
  assign _zz_5853 = _zz_5854;
  assign _zz_5854 = ($signed(data_mid_27_real) + $signed(_zz_573));
  assign _zz_5855 = _zz_5856;
  assign _zz_5856 = ($signed(_zz_5857) >>> _zz_576);
  assign _zz_5857 = _zz_5858;
  assign _zz_5858 = ($signed(data_mid_27_imag) + $signed(_zz_574));
  assign _zz_5859 = ($signed(twiddle_factor_table_3_real) * $signed(data_mid_36_real));
  assign _zz_5860 = ($signed(twiddle_factor_table_3_imag) * $signed(data_mid_36_imag));
  assign _zz_5861 = fixTo_288_dout;
  assign _zz_5862 = ($signed(twiddle_factor_table_3_real) * $signed(data_mid_36_imag));
  assign _zz_5863 = ($signed(twiddle_factor_table_3_imag) * $signed(data_mid_36_real));
  assign _zz_5864 = fixTo_289_dout;
  assign _zz_5865 = _zz_5866;
  assign _zz_5866 = ($signed(_zz_5867) >>> _zz_579);
  assign _zz_5867 = _zz_5868;
  assign _zz_5868 = ($signed(data_mid_32_real) - $signed(_zz_577));
  assign _zz_5869 = _zz_5870;
  assign _zz_5870 = ($signed(_zz_5871) >>> _zz_579);
  assign _zz_5871 = _zz_5872;
  assign _zz_5872 = ($signed(data_mid_32_imag) - $signed(_zz_578));
  assign _zz_5873 = _zz_5874;
  assign _zz_5874 = ($signed(_zz_5875) >>> _zz_580);
  assign _zz_5875 = _zz_5876;
  assign _zz_5876 = ($signed(data_mid_32_real) + $signed(_zz_577));
  assign _zz_5877 = _zz_5878;
  assign _zz_5878 = ($signed(_zz_5879) >>> _zz_580);
  assign _zz_5879 = _zz_5880;
  assign _zz_5880 = ($signed(data_mid_32_imag) + $signed(_zz_578));
  assign _zz_5881 = ($signed(twiddle_factor_table_4_real) * $signed(data_mid_37_real));
  assign _zz_5882 = ($signed(twiddle_factor_table_4_imag) * $signed(data_mid_37_imag));
  assign _zz_5883 = fixTo_290_dout;
  assign _zz_5884 = ($signed(twiddle_factor_table_4_real) * $signed(data_mid_37_imag));
  assign _zz_5885 = ($signed(twiddle_factor_table_4_imag) * $signed(data_mid_37_real));
  assign _zz_5886 = fixTo_291_dout;
  assign _zz_5887 = _zz_5888;
  assign _zz_5888 = ($signed(_zz_5889) >>> _zz_583);
  assign _zz_5889 = _zz_5890;
  assign _zz_5890 = ($signed(data_mid_33_real) - $signed(_zz_581));
  assign _zz_5891 = _zz_5892;
  assign _zz_5892 = ($signed(_zz_5893) >>> _zz_583);
  assign _zz_5893 = _zz_5894;
  assign _zz_5894 = ($signed(data_mid_33_imag) - $signed(_zz_582));
  assign _zz_5895 = _zz_5896;
  assign _zz_5896 = ($signed(_zz_5897) >>> _zz_584);
  assign _zz_5897 = _zz_5898;
  assign _zz_5898 = ($signed(data_mid_33_real) + $signed(_zz_581));
  assign _zz_5899 = _zz_5900;
  assign _zz_5900 = ($signed(_zz_5901) >>> _zz_584);
  assign _zz_5901 = _zz_5902;
  assign _zz_5902 = ($signed(data_mid_33_imag) + $signed(_zz_582));
  assign _zz_5903 = ($signed(twiddle_factor_table_5_real) * $signed(data_mid_38_real));
  assign _zz_5904 = ($signed(twiddle_factor_table_5_imag) * $signed(data_mid_38_imag));
  assign _zz_5905 = fixTo_292_dout;
  assign _zz_5906 = ($signed(twiddle_factor_table_5_real) * $signed(data_mid_38_imag));
  assign _zz_5907 = ($signed(twiddle_factor_table_5_imag) * $signed(data_mid_38_real));
  assign _zz_5908 = fixTo_293_dout;
  assign _zz_5909 = _zz_5910;
  assign _zz_5910 = ($signed(_zz_5911) >>> _zz_587);
  assign _zz_5911 = _zz_5912;
  assign _zz_5912 = ($signed(data_mid_34_real) - $signed(_zz_585));
  assign _zz_5913 = _zz_5914;
  assign _zz_5914 = ($signed(_zz_5915) >>> _zz_587);
  assign _zz_5915 = _zz_5916;
  assign _zz_5916 = ($signed(data_mid_34_imag) - $signed(_zz_586));
  assign _zz_5917 = _zz_5918;
  assign _zz_5918 = ($signed(_zz_5919) >>> _zz_588);
  assign _zz_5919 = _zz_5920;
  assign _zz_5920 = ($signed(data_mid_34_real) + $signed(_zz_585));
  assign _zz_5921 = _zz_5922;
  assign _zz_5922 = ($signed(_zz_5923) >>> _zz_588);
  assign _zz_5923 = _zz_5924;
  assign _zz_5924 = ($signed(data_mid_34_imag) + $signed(_zz_586));
  assign _zz_5925 = ($signed(twiddle_factor_table_6_real) * $signed(data_mid_39_real));
  assign _zz_5926 = ($signed(twiddle_factor_table_6_imag) * $signed(data_mid_39_imag));
  assign _zz_5927 = fixTo_294_dout;
  assign _zz_5928 = ($signed(twiddle_factor_table_6_real) * $signed(data_mid_39_imag));
  assign _zz_5929 = ($signed(twiddle_factor_table_6_imag) * $signed(data_mid_39_real));
  assign _zz_5930 = fixTo_295_dout;
  assign _zz_5931 = _zz_5932;
  assign _zz_5932 = ($signed(_zz_5933) >>> _zz_591);
  assign _zz_5933 = _zz_5934;
  assign _zz_5934 = ($signed(data_mid_35_real) - $signed(_zz_589));
  assign _zz_5935 = _zz_5936;
  assign _zz_5936 = ($signed(_zz_5937) >>> _zz_591);
  assign _zz_5937 = _zz_5938;
  assign _zz_5938 = ($signed(data_mid_35_imag) - $signed(_zz_590));
  assign _zz_5939 = _zz_5940;
  assign _zz_5940 = ($signed(_zz_5941) >>> _zz_592);
  assign _zz_5941 = _zz_5942;
  assign _zz_5942 = ($signed(data_mid_35_real) + $signed(_zz_589));
  assign _zz_5943 = _zz_5944;
  assign _zz_5944 = ($signed(_zz_5945) >>> _zz_592);
  assign _zz_5945 = _zz_5946;
  assign _zz_5946 = ($signed(data_mid_35_imag) + $signed(_zz_590));
  assign _zz_5947 = ($signed(twiddle_factor_table_3_real) * $signed(data_mid_44_real));
  assign _zz_5948 = ($signed(twiddle_factor_table_3_imag) * $signed(data_mid_44_imag));
  assign _zz_5949 = fixTo_296_dout;
  assign _zz_5950 = ($signed(twiddle_factor_table_3_real) * $signed(data_mid_44_imag));
  assign _zz_5951 = ($signed(twiddle_factor_table_3_imag) * $signed(data_mid_44_real));
  assign _zz_5952 = fixTo_297_dout;
  assign _zz_5953 = _zz_5954;
  assign _zz_5954 = ($signed(_zz_5955) >>> _zz_595);
  assign _zz_5955 = _zz_5956;
  assign _zz_5956 = ($signed(data_mid_40_real) - $signed(_zz_593));
  assign _zz_5957 = _zz_5958;
  assign _zz_5958 = ($signed(_zz_5959) >>> _zz_595);
  assign _zz_5959 = _zz_5960;
  assign _zz_5960 = ($signed(data_mid_40_imag) - $signed(_zz_594));
  assign _zz_5961 = _zz_5962;
  assign _zz_5962 = ($signed(_zz_5963) >>> _zz_596);
  assign _zz_5963 = _zz_5964;
  assign _zz_5964 = ($signed(data_mid_40_real) + $signed(_zz_593));
  assign _zz_5965 = _zz_5966;
  assign _zz_5966 = ($signed(_zz_5967) >>> _zz_596);
  assign _zz_5967 = _zz_5968;
  assign _zz_5968 = ($signed(data_mid_40_imag) + $signed(_zz_594));
  assign _zz_5969 = ($signed(twiddle_factor_table_4_real) * $signed(data_mid_45_real));
  assign _zz_5970 = ($signed(twiddle_factor_table_4_imag) * $signed(data_mid_45_imag));
  assign _zz_5971 = fixTo_298_dout;
  assign _zz_5972 = ($signed(twiddle_factor_table_4_real) * $signed(data_mid_45_imag));
  assign _zz_5973 = ($signed(twiddle_factor_table_4_imag) * $signed(data_mid_45_real));
  assign _zz_5974 = fixTo_299_dout;
  assign _zz_5975 = _zz_5976;
  assign _zz_5976 = ($signed(_zz_5977) >>> _zz_599);
  assign _zz_5977 = _zz_5978;
  assign _zz_5978 = ($signed(data_mid_41_real) - $signed(_zz_597));
  assign _zz_5979 = _zz_5980;
  assign _zz_5980 = ($signed(_zz_5981) >>> _zz_599);
  assign _zz_5981 = _zz_5982;
  assign _zz_5982 = ($signed(data_mid_41_imag) - $signed(_zz_598));
  assign _zz_5983 = _zz_5984;
  assign _zz_5984 = ($signed(_zz_5985) >>> _zz_600);
  assign _zz_5985 = _zz_5986;
  assign _zz_5986 = ($signed(data_mid_41_real) + $signed(_zz_597));
  assign _zz_5987 = _zz_5988;
  assign _zz_5988 = ($signed(_zz_5989) >>> _zz_600);
  assign _zz_5989 = _zz_5990;
  assign _zz_5990 = ($signed(data_mid_41_imag) + $signed(_zz_598));
  assign _zz_5991 = ($signed(twiddle_factor_table_5_real) * $signed(data_mid_46_real));
  assign _zz_5992 = ($signed(twiddle_factor_table_5_imag) * $signed(data_mid_46_imag));
  assign _zz_5993 = fixTo_300_dout;
  assign _zz_5994 = ($signed(twiddle_factor_table_5_real) * $signed(data_mid_46_imag));
  assign _zz_5995 = ($signed(twiddle_factor_table_5_imag) * $signed(data_mid_46_real));
  assign _zz_5996 = fixTo_301_dout;
  assign _zz_5997 = _zz_5998;
  assign _zz_5998 = ($signed(_zz_5999) >>> _zz_603);
  assign _zz_5999 = _zz_6000;
  assign _zz_6000 = ($signed(data_mid_42_real) - $signed(_zz_601));
  assign _zz_6001 = _zz_6002;
  assign _zz_6002 = ($signed(_zz_6003) >>> _zz_603);
  assign _zz_6003 = _zz_6004;
  assign _zz_6004 = ($signed(data_mid_42_imag) - $signed(_zz_602));
  assign _zz_6005 = _zz_6006;
  assign _zz_6006 = ($signed(_zz_6007) >>> _zz_604);
  assign _zz_6007 = _zz_6008;
  assign _zz_6008 = ($signed(data_mid_42_real) + $signed(_zz_601));
  assign _zz_6009 = _zz_6010;
  assign _zz_6010 = ($signed(_zz_6011) >>> _zz_604);
  assign _zz_6011 = _zz_6012;
  assign _zz_6012 = ($signed(data_mid_42_imag) + $signed(_zz_602));
  assign _zz_6013 = ($signed(twiddle_factor_table_6_real) * $signed(data_mid_47_real));
  assign _zz_6014 = ($signed(twiddle_factor_table_6_imag) * $signed(data_mid_47_imag));
  assign _zz_6015 = fixTo_302_dout;
  assign _zz_6016 = ($signed(twiddle_factor_table_6_real) * $signed(data_mid_47_imag));
  assign _zz_6017 = ($signed(twiddle_factor_table_6_imag) * $signed(data_mid_47_real));
  assign _zz_6018 = fixTo_303_dout;
  assign _zz_6019 = _zz_6020;
  assign _zz_6020 = ($signed(_zz_6021) >>> _zz_607);
  assign _zz_6021 = _zz_6022;
  assign _zz_6022 = ($signed(data_mid_43_real) - $signed(_zz_605));
  assign _zz_6023 = _zz_6024;
  assign _zz_6024 = ($signed(_zz_6025) >>> _zz_607);
  assign _zz_6025 = _zz_6026;
  assign _zz_6026 = ($signed(data_mid_43_imag) - $signed(_zz_606));
  assign _zz_6027 = _zz_6028;
  assign _zz_6028 = ($signed(_zz_6029) >>> _zz_608);
  assign _zz_6029 = _zz_6030;
  assign _zz_6030 = ($signed(data_mid_43_real) + $signed(_zz_605));
  assign _zz_6031 = _zz_6032;
  assign _zz_6032 = ($signed(_zz_6033) >>> _zz_608);
  assign _zz_6033 = _zz_6034;
  assign _zz_6034 = ($signed(data_mid_43_imag) + $signed(_zz_606));
  assign _zz_6035 = ($signed(twiddle_factor_table_3_real) * $signed(data_mid_52_real));
  assign _zz_6036 = ($signed(twiddle_factor_table_3_imag) * $signed(data_mid_52_imag));
  assign _zz_6037 = fixTo_304_dout;
  assign _zz_6038 = ($signed(twiddle_factor_table_3_real) * $signed(data_mid_52_imag));
  assign _zz_6039 = ($signed(twiddle_factor_table_3_imag) * $signed(data_mid_52_real));
  assign _zz_6040 = fixTo_305_dout;
  assign _zz_6041 = _zz_6042;
  assign _zz_6042 = ($signed(_zz_6043) >>> _zz_611);
  assign _zz_6043 = _zz_6044;
  assign _zz_6044 = ($signed(data_mid_48_real) - $signed(_zz_609));
  assign _zz_6045 = _zz_6046;
  assign _zz_6046 = ($signed(_zz_6047) >>> _zz_611);
  assign _zz_6047 = _zz_6048;
  assign _zz_6048 = ($signed(data_mid_48_imag) - $signed(_zz_610));
  assign _zz_6049 = _zz_6050;
  assign _zz_6050 = ($signed(_zz_6051) >>> _zz_612);
  assign _zz_6051 = _zz_6052;
  assign _zz_6052 = ($signed(data_mid_48_real) + $signed(_zz_609));
  assign _zz_6053 = _zz_6054;
  assign _zz_6054 = ($signed(_zz_6055) >>> _zz_612);
  assign _zz_6055 = _zz_6056;
  assign _zz_6056 = ($signed(data_mid_48_imag) + $signed(_zz_610));
  assign _zz_6057 = ($signed(twiddle_factor_table_4_real) * $signed(data_mid_53_real));
  assign _zz_6058 = ($signed(twiddle_factor_table_4_imag) * $signed(data_mid_53_imag));
  assign _zz_6059 = fixTo_306_dout;
  assign _zz_6060 = ($signed(twiddle_factor_table_4_real) * $signed(data_mid_53_imag));
  assign _zz_6061 = ($signed(twiddle_factor_table_4_imag) * $signed(data_mid_53_real));
  assign _zz_6062 = fixTo_307_dout;
  assign _zz_6063 = _zz_6064;
  assign _zz_6064 = ($signed(_zz_6065) >>> _zz_615);
  assign _zz_6065 = _zz_6066;
  assign _zz_6066 = ($signed(data_mid_49_real) - $signed(_zz_613));
  assign _zz_6067 = _zz_6068;
  assign _zz_6068 = ($signed(_zz_6069) >>> _zz_615);
  assign _zz_6069 = _zz_6070;
  assign _zz_6070 = ($signed(data_mid_49_imag) - $signed(_zz_614));
  assign _zz_6071 = _zz_6072;
  assign _zz_6072 = ($signed(_zz_6073) >>> _zz_616);
  assign _zz_6073 = _zz_6074;
  assign _zz_6074 = ($signed(data_mid_49_real) + $signed(_zz_613));
  assign _zz_6075 = _zz_6076;
  assign _zz_6076 = ($signed(_zz_6077) >>> _zz_616);
  assign _zz_6077 = _zz_6078;
  assign _zz_6078 = ($signed(data_mid_49_imag) + $signed(_zz_614));
  assign _zz_6079 = ($signed(twiddle_factor_table_5_real) * $signed(data_mid_54_real));
  assign _zz_6080 = ($signed(twiddle_factor_table_5_imag) * $signed(data_mid_54_imag));
  assign _zz_6081 = fixTo_308_dout;
  assign _zz_6082 = ($signed(twiddle_factor_table_5_real) * $signed(data_mid_54_imag));
  assign _zz_6083 = ($signed(twiddle_factor_table_5_imag) * $signed(data_mid_54_real));
  assign _zz_6084 = fixTo_309_dout;
  assign _zz_6085 = _zz_6086;
  assign _zz_6086 = ($signed(_zz_6087) >>> _zz_619);
  assign _zz_6087 = _zz_6088;
  assign _zz_6088 = ($signed(data_mid_50_real) - $signed(_zz_617));
  assign _zz_6089 = _zz_6090;
  assign _zz_6090 = ($signed(_zz_6091) >>> _zz_619);
  assign _zz_6091 = _zz_6092;
  assign _zz_6092 = ($signed(data_mid_50_imag) - $signed(_zz_618));
  assign _zz_6093 = _zz_6094;
  assign _zz_6094 = ($signed(_zz_6095) >>> _zz_620);
  assign _zz_6095 = _zz_6096;
  assign _zz_6096 = ($signed(data_mid_50_real) + $signed(_zz_617));
  assign _zz_6097 = _zz_6098;
  assign _zz_6098 = ($signed(_zz_6099) >>> _zz_620);
  assign _zz_6099 = _zz_6100;
  assign _zz_6100 = ($signed(data_mid_50_imag) + $signed(_zz_618));
  assign _zz_6101 = ($signed(twiddle_factor_table_6_real) * $signed(data_mid_55_real));
  assign _zz_6102 = ($signed(twiddle_factor_table_6_imag) * $signed(data_mid_55_imag));
  assign _zz_6103 = fixTo_310_dout;
  assign _zz_6104 = ($signed(twiddle_factor_table_6_real) * $signed(data_mid_55_imag));
  assign _zz_6105 = ($signed(twiddle_factor_table_6_imag) * $signed(data_mid_55_real));
  assign _zz_6106 = fixTo_311_dout;
  assign _zz_6107 = _zz_6108;
  assign _zz_6108 = ($signed(_zz_6109) >>> _zz_623);
  assign _zz_6109 = _zz_6110;
  assign _zz_6110 = ($signed(data_mid_51_real) - $signed(_zz_621));
  assign _zz_6111 = _zz_6112;
  assign _zz_6112 = ($signed(_zz_6113) >>> _zz_623);
  assign _zz_6113 = _zz_6114;
  assign _zz_6114 = ($signed(data_mid_51_imag) - $signed(_zz_622));
  assign _zz_6115 = _zz_6116;
  assign _zz_6116 = ($signed(_zz_6117) >>> _zz_624);
  assign _zz_6117 = _zz_6118;
  assign _zz_6118 = ($signed(data_mid_51_real) + $signed(_zz_621));
  assign _zz_6119 = _zz_6120;
  assign _zz_6120 = ($signed(_zz_6121) >>> _zz_624);
  assign _zz_6121 = _zz_6122;
  assign _zz_6122 = ($signed(data_mid_51_imag) + $signed(_zz_622));
  assign _zz_6123 = ($signed(twiddle_factor_table_3_real) * $signed(data_mid_60_real));
  assign _zz_6124 = ($signed(twiddle_factor_table_3_imag) * $signed(data_mid_60_imag));
  assign _zz_6125 = fixTo_312_dout;
  assign _zz_6126 = ($signed(twiddle_factor_table_3_real) * $signed(data_mid_60_imag));
  assign _zz_6127 = ($signed(twiddle_factor_table_3_imag) * $signed(data_mid_60_real));
  assign _zz_6128 = fixTo_313_dout;
  assign _zz_6129 = _zz_6130;
  assign _zz_6130 = ($signed(_zz_6131) >>> _zz_627);
  assign _zz_6131 = _zz_6132;
  assign _zz_6132 = ($signed(data_mid_56_real) - $signed(_zz_625));
  assign _zz_6133 = _zz_6134;
  assign _zz_6134 = ($signed(_zz_6135) >>> _zz_627);
  assign _zz_6135 = _zz_6136;
  assign _zz_6136 = ($signed(data_mid_56_imag) - $signed(_zz_626));
  assign _zz_6137 = _zz_6138;
  assign _zz_6138 = ($signed(_zz_6139) >>> _zz_628);
  assign _zz_6139 = _zz_6140;
  assign _zz_6140 = ($signed(data_mid_56_real) + $signed(_zz_625));
  assign _zz_6141 = _zz_6142;
  assign _zz_6142 = ($signed(_zz_6143) >>> _zz_628);
  assign _zz_6143 = _zz_6144;
  assign _zz_6144 = ($signed(data_mid_56_imag) + $signed(_zz_626));
  assign _zz_6145 = ($signed(twiddle_factor_table_4_real) * $signed(data_mid_61_real));
  assign _zz_6146 = ($signed(twiddle_factor_table_4_imag) * $signed(data_mid_61_imag));
  assign _zz_6147 = fixTo_314_dout;
  assign _zz_6148 = ($signed(twiddle_factor_table_4_real) * $signed(data_mid_61_imag));
  assign _zz_6149 = ($signed(twiddle_factor_table_4_imag) * $signed(data_mid_61_real));
  assign _zz_6150 = fixTo_315_dout;
  assign _zz_6151 = _zz_6152;
  assign _zz_6152 = ($signed(_zz_6153) >>> _zz_631);
  assign _zz_6153 = _zz_6154;
  assign _zz_6154 = ($signed(data_mid_57_real) - $signed(_zz_629));
  assign _zz_6155 = _zz_6156;
  assign _zz_6156 = ($signed(_zz_6157) >>> _zz_631);
  assign _zz_6157 = _zz_6158;
  assign _zz_6158 = ($signed(data_mid_57_imag) - $signed(_zz_630));
  assign _zz_6159 = _zz_6160;
  assign _zz_6160 = ($signed(_zz_6161) >>> _zz_632);
  assign _zz_6161 = _zz_6162;
  assign _zz_6162 = ($signed(data_mid_57_real) + $signed(_zz_629));
  assign _zz_6163 = _zz_6164;
  assign _zz_6164 = ($signed(_zz_6165) >>> _zz_632);
  assign _zz_6165 = _zz_6166;
  assign _zz_6166 = ($signed(data_mid_57_imag) + $signed(_zz_630));
  assign _zz_6167 = ($signed(twiddle_factor_table_5_real) * $signed(data_mid_62_real));
  assign _zz_6168 = ($signed(twiddle_factor_table_5_imag) * $signed(data_mid_62_imag));
  assign _zz_6169 = fixTo_316_dout;
  assign _zz_6170 = ($signed(twiddle_factor_table_5_real) * $signed(data_mid_62_imag));
  assign _zz_6171 = ($signed(twiddle_factor_table_5_imag) * $signed(data_mid_62_real));
  assign _zz_6172 = fixTo_317_dout;
  assign _zz_6173 = _zz_6174;
  assign _zz_6174 = ($signed(_zz_6175) >>> _zz_635);
  assign _zz_6175 = _zz_6176;
  assign _zz_6176 = ($signed(data_mid_58_real) - $signed(_zz_633));
  assign _zz_6177 = _zz_6178;
  assign _zz_6178 = ($signed(_zz_6179) >>> _zz_635);
  assign _zz_6179 = _zz_6180;
  assign _zz_6180 = ($signed(data_mid_58_imag) - $signed(_zz_634));
  assign _zz_6181 = _zz_6182;
  assign _zz_6182 = ($signed(_zz_6183) >>> _zz_636);
  assign _zz_6183 = _zz_6184;
  assign _zz_6184 = ($signed(data_mid_58_real) + $signed(_zz_633));
  assign _zz_6185 = _zz_6186;
  assign _zz_6186 = ($signed(_zz_6187) >>> _zz_636);
  assign _zz_6187 = _zz_6188;
  assign _zz_6188 = ($signed(data_mid_58_imag) + $signed(_zz_634));
  assign _zz_6189 = ($signed(twiddle_factor_table_6_real) * $signed(data_mid_63_real));
  assign _zz_6190 = ($signed(twiddle_factor_table_6_imag) * $signed(data_mid_63_imag));
  assign _zz_6191 = fixTo_318_dout;
  assign _zz_6192 = ($signed(twiddle_factor_table_6_real) * $signed(data_mid_63_imag));
  assign _zz_6193 = ($signed(twiddle_factor_table_6_imag) * $signed(data_mid_63_real));
  assign _zz_6194 = fixTo_319_dout;
  assign _zz_6195 = _zz_6196;
  assign _zz_6196 = ($signed(_zz_6197) >>> _zz_639);
  assign _zz_6197 = _zz_6198;
  assign _zz_6198 = ($signed(data_mid_59_real) - $signed(_zz_637));
  assign _zz_6199 = _zz_6200;
  assign _zz_6200 = ($signed(_zz_6201) >>> _zz_639);
  assign _zz_6201 = _zz_6202;
  assign _zz_6202 = ($signed(data_mid_59_imag) - $signed(_zz_638));
  assign _zz_6203 = _zz_6204;
  assign _zz_6204 = ($signed(_zz_6205) >>> _zz_640);
  assign _zz_6205 = _zz_6206;
  assign _zz_6206 = ($signed(data_mid_59_real) + $signed(_zz_637));
  assign _zz_6207 = _zz_6208;
  assign _zz_6208 = ($signed(_zz_6209) >>> _zz_640);
  assign _zz_6209 = _zz_6210;
  assign _zz_6210 = ($signed(data_mid_59_imag) + $signed(_zz_638));
  assign _zz_6211 = ($signed(twiddle_factor_table_3_real) * $signed(data_mid_68_real));
  assign _zz_6212 = ($signed(twiddle_factor_table_3_imag) * $signed(data_mid_68_imag));
  assign _zz_6213 = fixTo_320_dout;
  assign _zz_6214 = ($signed(twiddle_factor_table_3_real) * $signed(data_mid_68_imag));
  assign _zz_6215 = ($signed(twiddle_factor_table_3_imag) * $signed(data_mid_68_real));
  assign _zz_6216 = fixTo_321_dout;
  assign _zz_6217 = _zz_6218;
  assign _zz_6218 = ($signed(_zz_6219) >>> _zz_643);
  assign _zz_6219 = _zz_6220;
  assign _zz_6220 = ($signed(data_mid_64_real) - $signed(_zz_641));
  assign _zz_6221 = _zz_6222;
  assign _zz_6222 = ($signed(_zz_6223) >>> _zz_643);
  assign _zz_6223 = _zz_6224;
  assign _zz_6224 = ($signed(data_mid_64_imag) - $signed(_zz_642));
  assign _zz_6225 = _zz_6226;
  assign _zz_6226 = ($signed(_zz_6227) >>> _zz_644);
  assign _zz_6227 = _zz_6228;
  assign _zz_6228 = ($signed(data_mid_64_real) + $signed(_zz_641));
  assign _zz_6229 = _zz_6230;
  assign _zz_6230 = ($signed(_zz_6231) >>> _zz_644);
  assign _zz_6231 = _zz_6232;
  assign _zz_6232 = ($signed(data_mid_64_imag) + $signed(_zz_642));
  assign _zz_6233 = ($signed(twiddle_factor_table_4_real) * $signed(data_mid_69_real));
  assign _zz_6234 = ($signed(twiddle_factor_table_4_imag) * $signed(data_mid_69_imag));
  assign _zz_6235 = fixTo_322_dout;
  assign _zz_6236 = ($signed(twiddle_factor_table_4_real) * $signed(data_mid_69_imag));
  assign _zz_6237 = ($signed(twiddle_factor_table_4_imag) * $signed(data_mid_69_real));
  assign _zz_6238 = fixTo_323_dout;
  assign _zz_6239 = _zz_6240;
  assign _zz_6240 = ($signed(_zz_6241) >>> _zz_647);
  assign _zz_6241 = _zz_6242;
  assign _zz_6242 = ($signed(data_mid_65_real) - $signed(_zz_645));
  assign _zz_6243 = _zz_6244;
  assign _zz_6244 = ($signed(_zz_6245) >>> _zz_647);
  assign _zz_6245 = _zz_6246;
  assign _zz_6246 = ($signed(data_mid_65_imag) - $signed(_zz_646));
  assign _zz_6247 = _zz_6248;
  assign _zz_6248 = ($signed(_zz_6249) >>> _zz_648);
  assign _zz_6249 = _zz_6250;
  assign _zz_6250 = ($signed(data_mid_65_real) + $signed(_zz_645));
  assign _zz_6251 = _zz_6252;
  assign _zz_6252 = ($signed(_zz_6253) >>> _zz_648);
  assign _zz_6253 = _zz_6254;
  assign _zz_6254 = ($signed(data_mid_65_imag) + $signed(_zz_646));
  assign _zz_6255 = ($signed(twiddle_factor_table_5_real) * $signed(data_mid_70_real));
  assign _zz_6256 = ($signed(twiddle_factor_table_5_imag) * $signed(data_mid_70_imag));
  assign _zz_6257 = fixTo_324_dout;
  assign _zz_6258 = ($signed(twiddle_factor_table_5_real) * $signed(data_mid_70_imag));
  assign _zz_6259 = ($signed(twiddle_factor_table_5_imag) * $signed(data_mid_70_real));
  assign _zz_6260 = fixTo_325_dout;
  assign _zz_6261 = _zz_6262;
  assign _zz_6262 = ($signed(_zz_6263) >>> _zz_651);
  assign _zz_6263 = _zz_6264;
  assign _zz_6264 = ($signed(data_mid_66_real) - $signed(_zz_649));
  assign _zz_6265 = _zz_6266;
  assign _zz_6266 = ($signed(_zz_6267) >>> _zz_651);
  assign _zz_6267 = _zz_6268;
  assign _zz_6268 = ($signed(data_mid_66_imag) - $signed(_zz_650));
  assign _zz_6269 = _zz_6270;
  assign _zz_6270 = ($signed(_zz_6271) >>> _zz_652);
  assign _zz_6271 = _zz_6272;
  assign _zz_6272 = ($signed(data_mid_66_real) + $signed(_zz_649));
  assign _zz_6273 = _zz_6274;
  assign _zz_6274 = ($signed(_zz_6275) >>> _zz_652);
  assign _zz_6275 = _zz_6276;
  assign _zz_6276 = ($signed(data_mid_66_imag) + $signed(_zz_650));
  assign _zz_6277 = ($signed(twiddle_factor_table_6_real) * $signed(data_mid_71_real));
  assign _zz_6278 = ($signed(twiddle_factor_table_6_imag) * $signed(data_mid_71_imag));
  assign _zz_6279 = fixTo_326_dout;
  assign _zz_6280 = ($signed(twiddle_factor_table_6_real) * $signed(data_mid_71_imag));
  assign _zz_6281 = ($signed(twiddle_factor_table_6_imag) * $signed(data_mid_71_real));
  assign _zz_6282 = fixTo_327_dout;
  assign _zz_6283 = _zz_6284;
  assign _zz_6284 = ($signed(_zz_6285) >>> _zz_655);
  assign _zz_6285 = _zz_6286;
  assign _zz_6286 = ($signed(data_mid_67_real) - $signed(_zz_653));
  assign _zz_6287 = _zz_6288;
  assign _zz_6288 = ($signed(_zz_6289) >>> _zz_655);
  assign _zz_6289 = _zz_6290;
  assign _zz_6290 = ($signed(data_mid_67_imag) - $signed(_zz_654));
  assign _zz_6291 = _zz_6292;
  assign _zz_6292 = ($signed(_zz_6293) >>> _zz_656);
  assign _zz_6293 = _zz_6294;
  assign _zz_6294 = ($signed(data_mid_67_real) + $signed(_zz_653));
  assign _zz_6295 = _zz_6296;
  assign _zz_6296 = ($signed(_zz_6297) >>> _zz_656);
  assign _zz_6297 = _zz_6298;
  assign _zz_6298 = ($signed(data_mid_67_imag) + $signed(_zz_654));
  assign _zz_6299 = ($signed(twiddle_factor_table_3_real) * $signed(data_mid_76_real));
  assign _zz_6300 = ($signed(twiddle_factor_table_3_imag) * $signed(data_mid_76_imag));
  assign _zz_6301 = fixTo_328_dout;
  assign _zz_6302 = ($signed(twiddle_factor_table_3_real) * $signed(data_mid_76_imag));
  assign _zz_6303 = ($signed(twiddle_factor_table_3_imag) * $signed(data_mid_76_real));
  assign _zz_6304 = fixTo_329_dout;
  assign _zz_6305 = _zz_6306;
  assign _zz_6306 = ($signed(_zz_6307) >>> _zz_659);
  assign _zz_6307 = _zz_6308;
  assign _zz_6308 = ($signed(data_mid_72_real) - $signed(_zz_657));
  assign _zz_6309 = _zz_6310;
  assign _zz_6310 = ($signed(_zz_6311) >>> _zz_659);
  assign _zz_6311 = _zz_6312;
  assign _zz_6312 = ($signed(data_mid_72_imag) - $signed(_zz_658));
  assign _zz_6313 = _zz_6314;
  assign _zz_6314 = ($signed(_zz_6315) >>> _zz_660);
  assign _zz_6315 = _zz_6316;
  assign _zz_6316 = ($signed(data_mid_72_real) + $signed(_zz_657));
  assign _zz_6317 = _zz_6318;
  assign _zz_6318 = ($signed(_zz_6319) >>> _zz_660);
  assign _zz_6319 = _zz_6320;
  assign _zz_6320 = ($signed(data_mid_72_imag) + $signed(_zz_658));
  assign _zz_6321 = ($signed(twiddle_factor_table_4_real) * $signed(data_mid_77_real));
  assign _zz_6322 = ($signed(twiddle_factor_table_4_imag) * $signed(data_mid_77_imag));
  assign _zz_6323 = fixTo_330_dout;
  assign _zz_6324 = ($signed(twiddle_factor_table_4_real) * $signed(data_mid_77_imag));
  assign _zz_6325 = ($signed(twiddle_factor_table_4_imag) * $signed(data_mid_77_real));
  assign _zz_6326 = fixTo_331_dout;
  assign _zz_6327 = _zz_6328;
  assign _zz_6328 = ($signed(_zz_6329) >>> _zz_663);
  assign _zz_6329 = _zz_6330;
  assign _zz_6330 = ($signed(data_mid_73_real) - $signed(_zz_661));
  assign _zz_6331 = _zz_6332;
  assign _zz_6332 = ($signed(_zz_6333) >>> _zz_663);
  assign _zz_6333 = _zz_6334;
  assign _zz_6334 = ($signed(data_mid_73_imag) - $signed(_zz_662));
  assign _zz_6335 = _zz_6336;
  assign _zz_6336 = ($signed(_zz_6337) >>> _zz_664);
  assign _zz_6337 = _zz_6338;
  assign _zz_6338 = ($signed(data_mid_73_real) + $signed(_zz_661));
  assign _zz_6339 = _zz_6340;
  assign _zz_6340 = ($signed(_zz_6341) >>> _zz_664);
  assign _zz_6341 = _zz_6342;
  assign _zz_6342 = ($signed(data_mid_73_imag) + $signed(_zz_662));
  assign _zz_6343 = ($signed(twiddle_factor_table_5_real) * $signed(data_mid_78_real));
  assign _zz_6344 = ($signed(twiddle_factor_table_5_imag) * $signed(data_mid_78_imag));
  assign _zz_6345 = fixTo_332_dout;
  assign _zz_6346 = ($signed(twiddle_factor_table_5_real) * $signed(data_mid_78_imag));
  assign _zz_6347 = ($signed(twiddle_factor_table_5_imag) * $signed(data_mid_78_real));
  assign _zz_6348 = fixTo_333_dout;
  assign _zz_6349 = _zz_6350;
  assign _zz_6350 = ($signed(_zz_6351) >>> _zz_667);
  assign _zz_6351 = _zz_6352;
  assign _zz_6352 = ($signed(data_mid_74_real) - $signed(_zz_665));
  assign _zz_6353 = _zz_6354;
  assign _zz_6354 = ($signed(_zz_6355) >>> _zz_667);
  assign _zz_6355 = _zz_6356;
  assign _zz_6356 = ($signed(data_mid_74_imag) - $signed(_zz_666));
  assign _zz_6357 = _zz_6358;
  assign _zz_6358 = ($signed(_zz_6359) >>> _zz_668);
  assign _zz_6359 = _zz_6360;
  assign _zz_6360 = ($signed(data_mid_74_real) + $signed(_zz_665));
  assign _zz_6361 = _zz_6362;
  assign _zz_6362 = ($signed(_zz_6363) >>> _zz_668);
  assign _zz_6363 = _zz_6364;
  assign _zz_6364 = ($signed(data_mid_74_imag) + $signed(_zz_666));
  assign _zz_6365 = ($signed(twiddle_factor_table_6_real) * $signed(data_mid_79_real));
  assign _zz_6366 = ($signed(twiddle_factor_table_6_imag) * $signed(data_mid_79_imag));
  assign _zz_6367 = fixTo_334_dout;
  assign _zz_6368 = ($signed(twiddle_factor_table_6_real) * $signed(data_mid_79_imag));
  assign _zz_6369 = ($signed(twiddle_factor_table_6_imag) * $signed(data_mid_79_real));
  assign _zz_6370 = fixTo_335_dout;
  assign _zz_6371 = _zz_6372;
  assign _zz_6372 = ($signed(_zz_6373) >>> _zz_671);
  assign _zz_6373 = _zz_6374;
  assign _zz_6374 = ($signed(data_mid_75_real) - $signed(_zz_669));
  assign _zz_6375 = _zz_6376;
  assign _zz_6376 = ($signed(_zz_6377) >>> _zz_671);
  assign _zz_6377 = _zz_6378;
  assign _zz_6378 = ($signed(data_mid_75_imag) - $signed(_zz_670));
  assign _zz_6379 = _zz_6380;
  assign _zz_6380 = ($signed(_zz_6381) >>> _zz_672);
  assign _zz_6381 = _zz_6382;
  assign _zz_6382 = ($signed(data_mid_75_real) + $signed(_zz_669));
  assign _zz_6383 = _zz_6384;
  assign _zz_6384 = ($signed(_zz_6385) >>> _zz_672);
  assign _zz_6385 = _zz_6386;
  assign _zz_6386 = ($signed(data_mid_75_imag) + $signed(_zz_670));
  assign _zz_6387 = ($signed(twiddle_factor_table_3_real) * $signed(data_mid_84_real));
  assign _zz_6388 = ($signed(twiddle_factor_table_3_imag) * $signed(data_mid_84_imag));
  assign _zz_6389 = fixTo_336_dout;
  assign _zz_6390 = ($signed(twiddle_factor_table_3_real) * $signed(data_mid_84_imag));
  assign _zz_6391 = ($signed(twiddle_factor_table_3_imag) * $signed(data_mid_84_real));
  assign _zz_6392 = fixTo_337_dout;
  assign _zz_6393 = _zz_6394;
  assign _zz_6394 = ($signed(_zz_6395) >>> _zz_675);
  assign _zz_6395 = _zz_6396;
  assign _zz_6396 = ($signed(data_mid_80_real) - $signed(_zz_673));
  assign _zz_6397 = _zz_6398;
  assign _zz_6398 = ($signed(_zz_6399) >>> _zz_675);
  assign _zz_6399 = _zz_6400;
  assign _zz_6400 = ($signed(data_mid_80_imag) - $signed(_zz_674));
  assign _zz_6401 = _zz_6402;
  assign _zz_6402 = ($signed(_zz_6403) >>> _zz_676);
  assign _zz_6403 = _zz_6404;
  assign _zz_6404 = ($signed(data_mid_80_real) + $signed(_zz_673));
  assign _zz_6405 = _zz_6406;
  assign _zz_6406 = ($signed(_zz_6407) >>> _zz_676);
  assign _zz_6407 = _zz_6408;
  assign _zz_6408 = ($signed(data_mid_80_imag) + $signed(_zz_674));
  assign _zz_6409 = ($signed(twiddle_factor_table_4_real) * $signed(data_mid_85_real));
  assign _zz_6410 = ($signed(twiddle_factor_table_4_imag) * $signed(data_mid_85_imag));
  assign _zz_6411 = fixTo_338_dout;
  assign _zz_6412 = ($signed(twiddle_factor_table_4_real) * $signed(data_mid_85_imag));
  assign _zz_6413 = ($signed(twiddle_factor_table_4_imag) * $signed(data_mid_85_real));
  assign _zz_6414 = fixTo_339_dout;
  assign _zz_6415 = _zz_6416;
  assign _zz_6416 = ($signed(_zz_6417) >>> _zz_679);
  assign _zz_6417 = _zz_6418;
  assign _zz_6418 = ($signed(data_mid_81_real) - $signed(_zz_677));
  assign _zz_6419 = _zz_6420;
  assign _zz_6420 = ($signed(_zz_6421) >>> _zz_679);
  assign _zz_6421 = _zz_6422;
  assign _zz_6422 = ($signed(data_mid_81_imag) - $signed(_zz_678));
  assign _zz_6423 = _zz_6424;
  assign _zz_6424 = ($signed(_zz_6425) >>> _zz_680);
  assign _zz_6425 = _zz_6426;
  assign _zz_6426 = ($signed(data_mid_81_real) + $signed(_zz_677));
  assign _zz_6427 = _zz_6428;
  assign _zz_6428 = ($signed(_zz_6429) >>> _zz_680);
  assign _zz_6429 = _zz_6430;
  assign _zz_6430 = ($signed(data_mid_81_imag) + $signed(_zz_678));
  assign _zz_6431 = ($signed(twiddle_factor_table_5_real) * $signed(data_mid_86_real));
  assign _zz_6432 = ($signed(twiddle_factor_table_5_imag) * $signed(data_mid_86_imag));
  assign _zz_6433 = fixTo_340_dout;
  assign _zz_6434 = ($signed(twiddle_factor_table_5_real) * $signed(data_mid_86_imag));
  assign _zz_6435 = ($signed(twiddle_factor_table_5_imag) * $signed(data_mid_86_real));
  assign _zz_6436 = fixTo_341_dout;
  assign _zz_6437 = _zz_6438;
  assign _zz_6438 = ($signed(_zz_6439) >>> _zz_683);
  assign _zz_6439 = _zz_6440;
  assign _zz_6440 = ($signed(data_mid_82_real) - $signed(_zz_681));
  assign _zz_6441 = _zz_6442;
  assign _zz_6442 = ($signed(_zz_6443) >>> _zz_683);
  assign _zz_6443 = _zz_6444;
  assign _zz_6444 = ($signed(data_mid_82_imag) - $signed(_zz_682));
  assign _zz_6445 = _zz_6446;
  assign _zz_6446 = ($signed(_zz_6447) >>> _zz_684);
  assign _zz_6447 = _zz_6448;
  assign _zz_6448 = ($signed(data_mid_82_real) + $signed(_zz_681));
  assign _zz_6449 = _zz_6450;
  assign _zz_6450 = ($signed(_zz_6451) >>> _zz_684);
  assign _zz_6451 = _zz_6452;
  assign _zz_6452 = ($signed(data_mid_82_imag) + $signed(_zz_682));
  assign _zz_6453 = ($signed(twiddle_factor_table_6_real) * $signed(data_mid_87_real));
  assign _zz_6454 = ($signed(twiddle_factor_table_6_imag) * $signed(data_mid_87_imag));
  assign _zz_6455 = fixTo_342_dout;
  assign _zz_6456 = ($signed(twiddle_factor_table_6_real) * $signed(data_mid_87_imag));
  assign _zz_6457 = ($signed(twiddle_factor_table_6_imag) * $signed(data_mid_87_real));
  assign _zz_6458 = fixTo_343_dout;
  assign _zz_6459 = _zz_6460;
  assign _zz_6460 = ($signed(_zz_6461) >>> _zz_687);
  assign _zz_6461 = _zz_6462;
  assign _zz_6462 = ($signed(data_mid_83_real) - $signed(_zz_685));
  assign _zz_6463 = _zz_6464;
  assign _zz_6464 = ($signed(_zz_6465) >>> _zz_687);
  assign _zz_6465 = _zz_6466;
  assign _zz_6466 = ($signed(data_mid_83_imag) - $signed(_zz_686));
  assign _zz_6467 = _zz_6468;
  assign _zz_6468 = ($signed(_zz_6469) >>> _zz_688);
  assign _zz_6469 = _zz_6470;
  assign _zz_6470 = ($signed(data_mid_83_real) + $signed(_zz_685));
  assign _zz_6471 = _zz_6472;
  assign _zz_6472 = ($signed(_zz_6473) >>> _zz_688);
  assign _zz_6473 = _zz_6474;
  assign _zz_6474 = ($signed(data_mid_83_imag) + $signed(_zz_686));
  assign _zz_6475 = ($signed(twiddle_factor_table_3_real) * $signed(data_mid_92_real));
  assign _zz_6476 = ($signed(twiddle_factor_table_3_imag) * $signed(data_mid_92_imag));
  assign _zz_6477 = fixTo_344_dout;
  assign _zz_6478 = ($signed(twiddle_factor_table_3_real) * $signed(data_mid_92_imag));
  assign _zz_6479 = ($signed(twiddle_factor_table_3_imag) * $signed(data_mid_92_real));
  assign _zz_6480 = fixTo_345_dout;
  assign _zz_6481 = _zz_6482;
  assign _zz_6482 = ($signed(_zz_6483) >>> _zz_691);
  assign _zz_6483 = _zz_6484;
  assign _zz_6484 = ($signed(data_mid_88_real) - $signed(_zz_689));
  assign _zz_6485 = _zz_6486;
  assign _zz_6486 = ($signed(_zz_6487) >>> _zz_691);
  assign _zz_6487 = _zz_6488;
  assign _zz_6488 = ($signed(data_mid_88_imag) - $signed(_zz_690));
  assign _zz_6489 = _zz_6490;
  assign _zz_6490 = ($signed(_zz_6491) >>> _zz_692);
  assign _zz_6491 = _zz_6492;
  assign _zz_6492 = ($signed(data_mid_88_real) + $signed(_zz_689));
  assign _zz_6493 = _zz_6494;
  assign _zz_6494 = ($signed(_zz_6495) >>> _zz_692);
  assign _zz_6495 = _zz_6496;
  assign _zz_6496 = ($signed(data_mid_88_imag) + $signed(_zz_690));
  assign _zz_6497 = ($signed(twiddle_factor_table_4_real) * $signed(data_mid_93_real));
  assign _zz_6498 = ($signed(twiddle_factor_table_4_imag) * $signed(data_mid_93_imag));
  assign _zz_6499 = fixTo_346_dout;
  assign _zz_6500 = ($signed(twiddle_factor_table_4_real) * $signed(data_mid_93_imag));
  assign _zz_6501 = ($signed(twiddle_factor_table_4_imag) * $signed(data_mid_93_real));
  assign _zz_6502 = fixTo_347_dout;
  assign _zz_6503 = _zz_6504;
  assign _zz_6504 = ($signed(_zz_6505) >>> _zz_695);
  assign _zz_6505 = _zz_6506;
  assign _zz_6506 = ($signed(data_mid_89_real) - $signed(_zz_693));
  assign _zz_6507 = _zz_6508;
  assign _zz_6508 = ($signed(_zz_6509) >>> _zz_695);
  assign _zz_6509 = _zz_6510;
  assign _zz_6510 = ($signed(data_mid_89_imag) - $signed(_zz_694));
  assign _zz_6511 = _zz_6512;
  assign _zz_6512 = ($signed(_zz_6513) >>> _zz_696);
  assign _zz_6513 = _zz_6514;
  assign _zz_6514 = ($signed(data_mid_89_real) + $signed(_zz_693));
  assign _zz_6515 = _zz_6516;
  assign _zz_6516 = ($signed(_zz_6517) >>> _zz_696);
  assign _zz_6517 = _zz_6518;
  assign _zz_6518 = ($signed(data_mid_89_imag) + $signed(_zz_694));
  assign _zz_6519 = ($signed(twiddle_factor_table_5_real) * $signed(data_mid_94_real));
  assign _zz_6520 = ($signed(twiddle_factor_table_5_imag) * $signed(data_mid_94_imag));
  assign _zz_6521 = fixTo_348_dout;
  assign _zz_6522 = ($signed(twiddle_factor_table_5_real) * $signed(data_mid_94_imag));
  assign _zz_6523 = ($signed(twiddle_factor_table_5_imag) * $signed(data_mid_94_real));
  assign _zz_6524 = fixTo_349_dout;
  assign _zz_6525 = _zz_6526;
  assign _zz_6526 = ($signed(_zz_6527) >>> _zz_699);
  assign _zz_6527 = _zz_6528;
  assign _zz_6528 = ($signed(data_mid_90_real) - $signed(_zz_697));
  assign _zz_6529 = _zz_6530;
  assign _zz_6530 = ($signed(_zz_6531) >>> _zz_699);
  assign _zz_6531 = _zz_6532;
  assign _zz_6532 = ($signed(data_mid_90_imag) - $signed(_zz_698));
  assign _zz_6533 = _zz_6534;
  assign _zz_6534 = ($signed(_zz_6535) >>> _zz_700);
  assign _zz_6535 = _zz_6536;
  assign _zz_6536 = ($signed(data_mid_90_real) + $signed(_zz_697));
  assign _zz_6537 = _zz_6538;
  assign _zz_6538 = ($signed(_zz_6539) >>> _zz_700);
  assign _zz_6539 = _zz_6540;
  assign _zz_6540 = ($signed(data_mid_90_imag) + $signed(_zz_698));
  assign _zz_6541 = ($signed(twiddle_factor_table_6_real) * $signed(data_mid_95_real));
  assign _zz_6542 = ($signed(twiddle_factor_table_6_imag) * $signed(data_mid_95_imag));
  assign _zz_6543 = fixTo_350_dout;
  assign _zz_6544 = ($signed(twiddle_factor_table_6_real) * $signed(data_mid_95_imag));
  assign _zz_6545 = ($signed(twiddle_factor_table_6_imag) * $signed(data_mid_95_real));
  assign _zz_6546 = fixTo_351_dout;
  assign _zz_6547 = _zz_6548;
  assign _zz_6548 = ($signed(_zz_6549) >>> _zz_703);
  assign _zz_6549 = _zz_6550;
  assign _zz_6550 = ($signed(data_mid_91_real) - $signed(_zz_701));
  assign _zz_6551 = _zz_6552;
  assign _zz_6552 = ($signed(_zz_6553) >>> _zz_703);
  assign _zz_6553 = _zz_6554;
  assign _zz_6554 = ($signed(data_mid_91_imag) - $signed(_zz_702));
  assign _zz_6555 = _zz_6556;
  assign _zz_6556 = ($signed(_zz_6557) >>> _zz_704);
  assign _zz_6557 = _zz_6558;
  assign _zz_6558 = ($signed(data_mid_91_real) + $signed(_zz_701));
  assign _zz_6559 = _zz_6560;
  assign _zz_6560 = ($signed(_zz_6561) >>> _zz_704);
  assign _zz_6561 = _zz_6562;
  assign _zz_6562 = ($signed(data_mid_91_imag) + $signed(_zz_702));
  assign _zz_6563 = ($signed(twiddle_factor_table_3_real) * $signed(data_mid_100_real));
  assign _zz_6564 = ($signed(twiddle_factor_table_3_imag) * $signed(data_mid_100_imag));
  assign _zz_6565 = fixTo_352_dout;
  assign _zz_6566 = ($signed(twiddle_factor_table_3_real) * $signed(data_mid_100_imag));
  assign _zz_6567 = ($signed(twiddle_factor_table_3_imag) * $signed(data_mid_100_real));
  assign _zz_6568 = fixTo_353_dout;
  assign _zz_6569 = _zz_6570;
  assign _zz_6570 = ($signed(_zz_6571) >>> _zz_707);
  assign _zz_6571 = _zz_6572;
  assign _zz_6572 = ($signed(data_mid_96_real) - $signed(_zz_705));
  assign _zz_6573 = _zz_6574;
  assign _zz_6574 = ($signed(_zz_6575) >>> _zz_707);
  assign _zz_6575 = _zz_6576;
  assign _zz_6576 = ($signed(data_mid_96_imag) - $signed(_zz_706));
  assign _zz_6577 = _zz_6578;
  assign _zz_6578 = ($signed(_zz_6579) >>> _zz_708);
  assign _zz_6579 = _zz_6580;
  assign _zz_6580 = ($signed(data_mid_96_real) + $signed(_zz_705));
  assign _zz_6581 = _zz_6582;
  assign _zz_6582 = ($signed(_zz_6583) >>> _zz_708);
  assign _zz_6583 = _zz_6584;
  assign _zz_6584 = ($signed(data_mid_96_imag) + $signed(_zz_706));
  assign _zz_6585 = ($signed(twiddle_factor_table_4_real) * $signed(data_mid_101_real));
  assign _zz_6586 = ($signed(twiddle_factor_table_4_imag) * $signed(data_mid_101_imag));
  assign _zz_6587 = fixTo_354_dout;
  assign _zz_6588 = ($signed(twiddle_factor_table_4_real) * $signed(data_mid_101_imag));
  assign _zz_6589 = ($signed(twiddle_factor_table_4_imag) * $signed(data_mid_101_real));
  assign _zz_6590 = fixTo_355_dout;
  assign _zz_6591 = _zz_6592;
  assign _zz_6592 = ($signed(_zz_6593) >>> _zz_711);
  assign _zz_6593 = _zz_6594;
  assign _zz_6594 = ($signed(data_mid_97_real) - $signed(_zz_709));
  assign _zz_6595 = _zz_6596;
  assign _zz_6596 = ($signed(_zz_6597) >>> _zz_711);
  assign _zz_6597 = _zz_6598;
  assign _zz_6598 = ($signed(data_mid_97_imag) - $signed(_zz_710));
  assign _zz_6599 = _zz_6600;
  assign _zz_6600 = ($signed(_zz_6601) >>> _zz_712);
  assign _zz_6601 = _zz_6602;
  assign _zz_6602 = ($signed(data_mid_97_real) + $signed(_zz_709));
  assign _zz_6603 = _zz_6604;
  assign _zz_6604 = ($signed(_zz_6605) >>> _zz_712);
  assign _zz_6605 = _zz_6606;
  assign _zz_6606 = ($signed(data_mid_97_imag) + $signed(_zz_710));
  assign _zz_6607 = ($signed(twiddle_factor_table_5_real) * $signed(data_mid_102_real));
  assign _zz_6608 = ($signed(twiddle_factor_table_5_imag) * $signed(data_mid_102_imag));
  assign _zz_6609 = fixTo_356_dout;
  assign _zz_6610 = ($signed(twiddle_factor_table_5_real) * $signed(data_mid_102_imag));
  assign _zz_6611 = ($signed(twiddle_factor_table_5_imag) * $signed(data_mid_102_real));
  assign _zz_6612 = fixTo_357_dout;
  assign _zz_6613 = _zz_6614;
  assign _zz_6614 = ($signed(_zz_6615) >>> _zz_715);
  assign _zz_6615 = _zz_6616;
  assign _zz_6616 = ($signed(data_mid_98_real) - $signed(_zz_713));
  assign _zz_6617 = _zz_6618;
  assign _zz_6618 = ($signed(_zz_6619) >>> _zz_715);
  assign _zz_6619 = _zz_6620;
  assign _zz_6620 = ($signed(data_mid_98_imag) - $signed(_zz_714));
  assign _zz_6621 = _zz_6622;
  assign _zz_6622 = ($signed(_zz_6623) >>> _zz_716);
  assign _zz_6623 = _zz_6624;
  assign _zz_6624 = ($signed(data_mid_98_real) + $signed(_zz_713));
  assign _zz_6625 = _zz_6626;
  assign _zz_6626 = ($signed(_zz_6627) >>> _zz_716);
  assign _zz_6627 = _zz_6628;
  assign _zz_6628 = ($signed(data_mid_98_imag) + $signed(_zz_714));
  assign _zz_6629 = ($signed(twiddle_factor_table_6_real) * $signed(data_mid_103_real));
  assign _zz_6630 = ($signed(twiddle_factor_table_6_imag) * $signed(data_mid_103_imag));
  assign _zz_6631 = fixTo_358_dout;
  assign _zz_6632 = ($signed(twiddle_factor_table_6_real) * $signed(data_mid_103_imag));
  assign _zz_6633 = ($signed(twiddle_factor_table_6_imag) * $signed(data_mid_103_real));
  assign _zz_6634 = fixTo_359_dout;
  assign _zz_6635 = _zz_6636;
  assign _zz_6636 = ($signed(_zz_6637) >>> _zz_719);
  assign _zz_6637 = _zz_6638;
  assign _zz_6638 = ($signed(data_mid_99_real) - $signed(_zz_717));
  assign _zz_6639 = _zz_6640;
  assign _zz_6640 = ($signed(_zz_6641) >>> _zz_719);
  assign _zz_6641 = _zz_6642;
  assign _zz_6642 = ($signed(data_mid_99_imag) - $signed(_zz_718));
  assign _zz_6643 = _zz_6644;
  assign _zz_6644 = ($signed(_zz_6645) >>> _zz_720);
  assign _zz_6645 = _zz_6646;
  assign _zz_6646 = ($signed(data_mid_99_real) + $signed(_zz_717));
  assign _zz_6647 = _zz_6648;
  assign _zz_6648 = ($signed(_zz_6649) >>> _zz_720);
  assign _zz_6649 = _zz_6650;
  assign _zz_6650 = ($signed(data_mid_99_imag) + $signed(_zz_718));
  assign _zz_6651 = ($signed(twiddle_factor_table_3_real) * $signed(data_mid_108_real));
  assign _zz_6652 = ($signed(twiddle_factor_table_3_imag) * $signed(data_mid_108_imag));
  assign _zz_6653 = fixTo_360_dout;
  assign _zz_6654 = ($signed(twiddle_factor_table_3_real) * $signed(data_mid_108_imag));
  assign _zz_6655 = ($signed(twiddle_factor_table_3_imag) * $signed(data_mid_108_real));
  assign _zz_6656 = fixTo_361_dout;
  assign _zz_6657 = _zz_6658;
  assign _zz_6658 = ($signed(_zz_6659) >>> _zz_723);
  assign _zz_6659 = _zz_6660;
  assign _zz_6660 = ($signed(data_mid_104_real) - $signed(_zz_721));
  assign _zz_6661 = _zz_6662;
  assign _zz_6662 = ($signed(_zz_6663) >>> _zz_723);
  assign _zz_6663 = _zz_6664;
  assign _zz_6664 = ($signed(data_mid_104_imag) - $signed(_zz_722));
  assign _zz_6665 = _zz_6666;
  assign _zz_6666 = ($signed(_zz_6667) >>> _zz_724);
  assign _zz_6667 = _zz_6668;
  assign _zz_6668 = ($signed(data_mid_104_real) + $signed(_zz_721));
  assign _zz_6669 = _zz_6670;
  assign _zz_6670 = ($signed(_zz_6671) >>> _zz_724);
  assign _zz_6671 = _zz_6672;
  assign _zz_6672 = ($signed(data_mid_104_imag) + $signed(_zz_722));
  assign _zz_6673 = ($signed(twiddle_factor_table_4_real) * $signed(data_mid_109_real));
  assign _zz_6674 = ($signed(twiddle_factor_table_4_imag) * $signed(data_mid_109_imag));
  assign _zz_6675 = fixTo_362_dout;
  assign _zz_6676 = ($signed(twiddle_factor_table_4_real) * $signed(data_mid_109_imag));
  assign _zz_6677 = ($signed(twiddle_factor_table_4_imag) * $signed(data_mid_109_real));
  assign _zz_6678 = fixTo_363_dout;
  assign _zz_6679 = _zz_6680;
  assign _zz_6680 = ($signed(_zz_6681) >>> _zz_727);
  assign _zz_6681 = _zz_6682;
  assign _zz_6682 = ($signed(data_mid_105_real) - $signed(_zz_725));
  assign _zz_6683 = _zz_6684;
  assign _zz_6684 = ($signed(_zz_6685) >>> _zz_727);
  assign _zz_6685 = _zz_6686;
  assign _zz_6686 = ($signed(data_mid_105_imag) - $signed(_zz_726));
  assign _zz_6687 = _zz_6688;
  assign _zz_6688 = ($signed(_zz_6689) >>> _zz_728);
  assign _zz_6689 = _zz_6690;
  assign _zz_6690 = ($signed(data_mid_105_real) + $signed(_zz_725));
  assign _zz_6691 = _zz_6692;
  assign _zz_6692 = ($signed(_zz_6693) >>> _zz_728);
  assign _zz_6693 = _zz_6694;
  assign _zz_6694 = ($signed(data_mid_105_imag) + $signed(_zz_726));
  assign _zz_6695 = ($signed(twiddle_factor_table_5_real) * $signed(data_mid_110_real));
  assign _zz_6696 = ($signed(twiddle_factor_table_5_imag) * $signed(data_mid_110_imag));
  assign _zz_6697 = fixTo_364_dout;
  assign _zz_6698 = ($signed(twiddle_factor_table_5_real) * $signed(data_mid_110_imag));
  assign _zz_6699 = ($signed(twiddle_factor_table_5_imag) * $signed(data_mid_110_real));
  assign _zz_6700 = fixTo_365_dout;
  assign _zz_6701 = _zz_6702;
  assign _zz_6702 = ($signed(_zz_6703) >>> _zz_731);
  assign _zz_6703 = _zz_6704;
  assign _zz_6704 = ($signed(data_mid_106_real) - $signed(_zz_729));
  assign _zz_6705 = _zz_6706;
  assign _zz_6706 = ($signed(_zz_6707) >>> _zz_731);
  assign _zz_6707 = _zz_6708;
  assign _zz_6708 = ($signed(data_mid_106_imag) - $signed(_zz_730));
  assign _zz_6709 = _zz_6710;
  assign _zz_6710 = ($signed(_zz_6711) >>> _zz_732);
  assign _zz_6711 = _zz_6712;
  assign _zz_6712 = ($signed(data_mid_106_real) + $signed(_zz_729));
  assign _zz_6713 = _zz_6714;
  assign _zz_6714 = ($signed(_zz_6715) >>> _zz_732);
  assign _zz_6715 = _zz_6716;
  assign _zz_6716 = ($signed(data_mid_106_imag) + $signed(_zz_730));
  assign _zz_6717 = ($signed(twiddle_factor_table_6_real) * $signed(data_mid_111_real));
  assign _zz_6718 = ($signed(twiddle_factor_table_6_imag) * $signed(data_mid_111_imag));
  assign _zz_6719 = fixTo_366_dout;
  assign _zz_6720 = ($signed(twiddle_factor_table_6_real) * $signed(data_mid_111_imag));
  assign _zz_6721 = ($signed(twiddle_factor_table_6_imag) * $signed(data_mid_111_real));
  assign _zz_6722 = fixTo_367_dout;
  assign _zz_6723 = _zz_6724;
  assign _zz_6724 = ($signed(_zz_6725) >>> _zz_735);
  assign _zz_6725 = _zz_6726;
  assign _zz_6726 = ($signed(data_mid_107_real) - $signed(_zz_733));
  assign _zz_6727 = _zz_6728;
  assign _zz_6728 = ($signed(_zz_6729) >>> _zz_735);
  assign _zz_6729 = _zz_6730;
  assign _zz_6730 = ($signed(data_mid_107_imag) - $signed(_zz_734));
  assign _zz_6731 = _zz_6732;
  assign _zz_6732 = ($signed(_zz_6733) >>> _zz_736);
  assign _zz_6733 = _zz_6734;
  assign _zz_6734 = ($signed(data_mid_107_real) + $signed(_zz_733));
  assign _zz_6735 = _zz_6736;
  assign _zz_6736 = ($signed(_zz_6737) >>> _zz_736);
  assign _zz_6737 = _zz_6738;
  assign _zz_6738 = ($signed(data_mid_107_imag) + $signed(_zz_734));
  assign _zz_6739 = ($signed(twiddle_factor_table_3_real) * $signed(data_mid_116_real));
  assign _zz_6740 = ($signed(twiddle_factor_table_3_imag) * $signed(data_mid_116_imag));
  assign _zz_6741 = fixTo_368_dout;
  assign _zz_6742 = ($signed(twiddle_factor_table_3_real) * $signed(data_mid_116_imag));
  assign _zz_6743 = ($signed(twiddle_factor_table_3_imag) * $signed(data_mid_116_real));
  assign _zz_6744 = fixTo_369_dout;
  assign _zz_6745 = _zz_6746;
  assign _zz_6746 = ($signed(_zz_6747) >>> _zz_739);
  assign _zz_6747 = _zz_6748;
  assign _zz_6748 = ($signed(data_mid_112_real) - $signed(_zz_737));
  assign _zz_6749 = _zz_6750;
  assign _zz_6750 = ($signed(_zz_6751) >>> _zz_739);
  assign _zz_6751 = _zz_6752;
  assign _zz_6752 = ($signed(data_mid_112_imag) - $signed(_zz_738));
  assign _zz_6753 = _zz_6754;
  assign _zz_6754 = ($signed(_zz_6755) >>> _zz_740);
  assign _zz_6755 = _zz_6756;
  assign _zz_6756 = ($signed(data_mid_112_real) + $signed(_zz_737));
  assign _zz_6757 = _zz_6758;
  assign _zz_6758 = ($signed(_zz_6759) >>> _zz_740);
  assign _zz_6759 = _zz_6760;
  assign _zz_6760 = ($signed(data_mid_112_imag) + $signed(_zz_738));
  assign _zz_6761 = ($signed(twiddle_factor_table_4_real) * $signed(data_mid_117_real));
  assign _zz_6762 = ($signed(twiddle_factor_table_4_imag) * $signed(data_mid_117_imag));
  assign _zz_6763 = fixTo_370_dout;
  assign _zz_6764 = ($signed(twiddle_factor_table_4_real) * $signed(data_mid_117_imag));
  assign _zz_6765 = ($signed(twiddle_factor_table_4_imag) * $signed(data_mid_117_real));
  assign _zz_6766 = fixTo_371_dout;
  assign _zz_6767 = _zz_6768;
  assign _zz_6768 = ($signed(_zz_6769) >>> _zz_743);
  assign _zz_6769 = _zz_6770;
  assign _zz_6770 = ($signed(data_mid_113_real) - $signed(_zz_741));
  assign _zz_6771 = _zz_6772;
  assign _zz_6772 = ($signed(_zz_6773) >>> _zz_743);
  assign _zz_6773 = _zz_6774;
  assign _zz_6774 = ($signed(data_mid_113_imag) - $signed(_zz_742));
  assign _zz_6775 = _zz_6776;
  assign _zz_6776 = ($signed(_zz_6777) >>> _zz_744);
  assign _zz_6777 = _zz_6778;
  assign _zz_6778 = ($signed(data_mid_113_real) + $signed(_zz_741));
  assign _zz_6779 = _zz_6780;
  assign _zz_6780 = ($signed(_zz_6781) >>> _zz_744);
  assign _zz_6781 = _zz_6782;
  assign _zz_6782 = ($signed(data_mid_113_imag) + $signed(_zz_742));
  assign _zz_6783 = ($signed(twiddle_factor_table_5_real) * $signed(data_mid_118_real));
  assign _zz_6784 = ($signed(twiddle_factor_table_5_imag) * $signed(data_mid_118_imag));
  assign _zz_6785 = fixTo_372_dout;
  assign _zz_6786 = ($signed(twiddle_factor_table_5_real) * $signed(data_mid_118_imag));
  assign _zz_6787 = ($signed(twiddle_factor_table_5_imag) * $signed(data_mid_118_real));
  assign _zz_6788 = fixTo_373_dout;
  assign _zz_6789 = _zz_6790;
  assign _zz_6790 = ($signed(_zz_6791) >>> _zz_747);
  assign _zz_6791 = _zz_6792;
  assign _zz_6792 = ($signed(data_mid_114_real) - $signed(_zz_745));
  assign _zz_6793 = _zz_6794;
  assign _zz_6794 = ($signed(_zz_6795) >>> _zz_747);
  assign _zz_6795 = _zz_6796;
  assign _zz_6796 = ($signed(data_mid_114_imag) - $signed(_zz_746));
  assign _zz_6797 = _zz_6798;
  assign _zz_6798 = ($signed(_zz_6799) >>> _zz_748);
  assign _zz_6799 = _zz_6800;
  assign _zz_6800 = ($signed(data_mid_114_real) + $signed(_zz_745));
  assign _zz_6801 = _zz_6802;
  assign _zz_6802 = ($signed(_zz_6803) >>> _zz_748);
  assign _zz_6803 = _zz_6804;
  assign _zz_6804 = ($signed(data_mid_114_imag) + $signed(_zz_746));
  assign _zz_6805 = ($signed(twiddle_factor_table_6_real) * $signed(data_mid_119_real));
  assign _zz_6806 = ($signed(twiddle_factor_table_6_imag) * $signed(data_mid_119_imag));
  assign _zz_6807 = fixTo_374_dout;
  assign _zz_6808 = ($signed(twiddle_factor_table_6_real) * $signed(data_mid_119_imag));
  assign _zz_6809 = ($signed(twiddle_factor_table_6_imag) * $signed(data_mid_119_real));
  assign _zz_6810 = fixTo_375_dout;
  assign _zz_6811 = _zz_6812;
  assign _zz_6812 = ($signed(_zz_6813) >>> _zz_751);
  assign _zz_6813 = _zz_6814;
  assign _zz_6814 = ($signed(data_mid_115_real) - $signed(_zz_749));
  assign _zz_6815 = _zz_6816;
  assign _zz_6816 = ($signed(_zz_6817) >>> _zz_751);
  assign _zz_6817 = _zz_6818;
  assign _zz_6818 = ($signed(data_mid_115_imag) - $signed(_zz_750));
  assign _zz_6819 = _zz_6820;
  assign _zz_6820 = ($signed(_zz_6821) >>> _zz_752);
  assign _zz_6821 = _zz_6822;
  assign _zz_6822 = ($signed(data_mid_115_real) + $signed(_zz_749));
  assign _zz_6823 = _zz_6824;
  assign _zz_6824 = ($signed(_zz_6825) >>> _zz_752);
  assign _zz_6825 = _zz_6826;
  assign _zz_6826 = ($signed(data_mid_115_imag) + $signed(_zz_750));
  assign _zz_6827 = ($signed(twiddle_factor_table_3_real) * $signed(data_mid_124_real));
  assign _zz_6828 = ($signed(twiddle_factor_table_3_imag) * $signed(data_mid_124_imag));
  assign _zz_6829 = fixTo_376_dout;
  assign _zz_6830 = ($signed(twiddle_factor_table_3_real) * $signed(data_mid_124_imag));
  assign _zz_6831 = ($signed(twiddle_factor_table_3_imag) * $signed(data_mid_124_real));
  assign _zz_6832 = fixTo_377_dout;
  assign _zz_6833 = _zz_6834;
  assign _zz_6834 = ($signed(_zz_6835) >>> _zz_755);
  assign _zz_6835 = _zz_6836;
  assign _zz_6836 = ($signed(data_mid_120_real) - $signed(_zz_753));
  assign _zz_6837 = _zz_6838;
  assign _zz_6838 = ($signed(_zz_6839) >>> _zz_755);
  assign _zz_6839 = _zz_6840;
  assign _zz_6840 = ($signed(data_mid_120_imag) - $signed(_zz_754));
  assign _zz_6841 = _zz_6842;
  assign _zz_6842 = ($signed(_zz_6843) >>> _zz_756);
  assign _zz_6843 = _zz_6844;
  assign _zz_6844 = ($signed(data_mid_120_real) + $signed(_zz_753));
  assign _zz_6845 = _zz_6846;
  assign _zz_6846 = ($signed(_zz_6847) >>> _zz_756);
  assign _zz_6847 = _zz_6848;
  assign _zz_6848 = ($signed(data_mid_120_imag) + $signed(_zz_754));
  assign _zz_6849 = ($signed(twiddle_factor_table_4_real) * $signed(data_mid_125_real));
  assign _zz_6850 = ($signed(twiddle_factor_table_4_imag) * $signed(data_mid_125_imag));
  assign _zz_6851 = fixTo_378_dout;
  assign _zz_6852 = ($signed(twiddle_factor_table_4_real) * $signed(data_mid_125_imag));
  assign _zz_6853 = ($signed(twiddle_factor_table_4_imag) * $signed(data_mid_125_real));
  assign _zz_6854 = fixTo_379_dout;
  assign _zz_6855 = _zz_6856;
  assign _zz_6856 = ($signed(_zz_6857) >>> _zz_759);
  assign _zz_6857 = _zz_6858;
  assign _zz_6858 = ($signed(data_mid_121_real) - $signed(_zz_757));
  assign _zz_6859 = _zz_6860;
  assign _zz_6860 = ($signed(_zz_6861) >>> _zz_759);
  assign _zz_6861 = _zz_6862;
  assign _zz_6862 = ($signed(data_mid_121_imag) - $signed(_zz_758));
  assign _zz_6863 = _zz_6864;
  assign _zz_6864 = ($signed(_zz_6865) >>> _zz_760);
  assign _zz_6865 = _zz_6866;
  assign _zz_6866 = ($signed(data_mid_121_real) + $signed(_zz_757));
  assign _zz_6867 = _zz_6868;
  assign _zz_6868 = ($signed(_zz_6869) >>> _zz_760);
  assign _zz_6869 = _zz_6870;
  assign _zz_6870 = ($signed(data_mid_121_imag) + $signed(_zz_758));
  assign _zz_6871 = ($signed(twiddle_factor_table_5_real) * $signed(data_mid_126_real));
  assign _zz_6872 = ($signed(twiddle_factor_table_5_imag) * $signed(data_mid_126_imag));
  assign _zz_6873 = fixTo_380_dout;
  assign _zz_6874 = ($signed(twiddle_factor_table_5_real) * $signed(data_mid_126_imag));
  assign _zz_6875 = ($signed(twiddle_factor_table_5_imag) * $signed(data_mid_126_real));
  assign _zz_6876 = fixTo_381_dout;
  assign _zz_6877 = _zz_6878;
  assign _zz_6878 = ($signed(_zz_6879) >>> _zz_763);
  assign _zz_6879 = _zz_6880;
  assign _zz_6880 = ($signed(data_mid_122_real) - $signed(_zz_761));
  assign _zz_6881 = _zz_6882;
  assign _zz_6882 = ($signed(_zz_6883) >>> _zz_763);
  assign _zz_6883 = _zz_6884;
  assign _zz_6884 = ($signed(data_mid_122_imag) - $signed(_zz_762));
  assign _zz_6885 = _zz_6886;
  assign _zz_6886 = ($signed(_zz_6887) >>> _zz_764);
  assign _zz_6887 = _zz_6888;
  assign _zz_6888 = ($signed(data_mid_122_real) + $signed(_zz_761));
  assign _zz_6889 = _zz_6890;
  assign _zz_6890 = ($signed(_zz_6891) >>> _zz_764);
  assign _zz_6891 = _zz_6892;
  assign _zz_6892 = ($signed(data_mid_122_imag) + $signed(_zz_762));
  assign _zz_6893 = ($signed(twiddle_factor_table_6_real) * $signed(data_mid_127_real));
  assign _zz_6894 = ($signed(twiddle_factor_table_6_imag) * $signed(data_mid_127_imag));
  assign _zz_6895 = fixTo_382_dout;
  assign _zz_6896 = ($signed(twiddle_factor_table_6_real) * $signed(data_mid_127_imag));
  assign _zz_6897 = ($signed(twiddle_factor_table_6_imag) * $signed(data_mid_127_real));
  assign _zz_6898 = fixTo_383_dout;
  assign _zz_6899 = _zz_6900;
  assign _zz_6900 = ($signed(_zz_6901) >>> _zz_767);
  assign _zz_6901 = _zz_6902;
  assign _zz_6902 = ($signed(data_mid_123_real) - $signed(_zz_765));
  assign _zz_6903 = _zz_6904;
  assign _zz_6904 = ($signed(_zz_6905) >>> _zz_767);
  assign _zz_6905 = _zz_6906;
  assign _zz_6906 = ($signed(data_mid_123_imag) - $signed(_zz_766));
  assign _zz_6907 = _zz_6908;
  assign _zz_6908 = ($signed(_zz_6909) >>> _zz_768);
  assign _zz_6909 = _zz_6910;
  assign _zz_6910 = ($signed(data_mid_123_real) + $signed(_zz_765));
  assign _zz_6911 = _zz_6912;
  assign _zz_6912 = ($signed(_zz_6913) >>> _zz_768);
  assign _zz_6913 = _zz_6914;
  assign _zz_6914 = ($signed(data_mid_123_imag) + $signed(_zz_766));
  assign _zz_6915 = ($signed(twiddle_factor_table_7_real) * $signed(data_mid_8_real));
  assign _zz_6916 = ($signed(twiddle_factor_table_7_imag) * $signed(data_mid_8_imag));
  assign _zz_6917 = fixTo_384_dout;
  assign _zz_6918 = ($signed(twiddle_factor_table_7_real) * $signed(data_mid_8_imag));
  assign _zz_6919 = ($signed(twiddle_factor_table_7_imag) * $signed(data_mid_8_real));
  assign _zz_6920 = fixTo_385_dout;
  assign _zz_6921 = _zz_6922;
  assign _zz_6922 = ($signed(_zz_6923) >>> _zz_771);
  assign _zz_6923 = _zz_6924;
  assign _zz_6924 = ($signed(data_mid_0_real) - $signed(_zz_769));
  assign _zz_6925 = _zz_6926;
  assign _zz_6926 = ($signed(_zz_6927) >>> _zz_771);
  assign _zz_6927 = _zz_6928;
  assign _zz_6928 = ($signed(data_mid_0_imag) - $signed(_zz_770));
  assign _zz_6929 = _zz_6930;
  assign _zz_6930 = ($signed(_zz_6931) >>> _zz_772);
  assign _zz_6931 = _zz_6932;
  assign _zz_6932 = ($signed(data_mid_0_real) + $signed(_zz_769));
  assign _zz_6933 = _zz_6934;
  assign _zz_6934 = ($signed(_zz_6935) >>> _zz_772);
  assign _zz_6935 = _zz_6936;
  assign _zz_6936 = ($signed(data_mid_0_imag) + $signed(_zz_770));
  assign _zz_6937 = ($signed(twiddle_factor_table_8_real) * $signed(data_mid_9_real));
  assign _zz_6938 = ($signed(twiddle_factor_table_8_imag) * $signed(data_mid_9_imag));
  assign _zz_6939 = fixTo_386_dout;
  assign _zz_6940 = ($signed(twiddle_factor_table_8_real) * $signed(data_mid_9_imag));
  assign _zz_6941 = ($signed(twiddle_factor_table_8_imag) * $signed(data_mid_9_real));
  assign _zz_6942 = fixTo_387_dout;
  assign _zz_6943 = _zz_6944;
  assign _zz_6944 = ($signed(_zz_6945) >>> _zz_775);
  assign _zz_6945 = _zz_6946;
  assign _zz_6946 = ($signed(data_mid_1_real) - $signed(_zz_773));
  assign _zz_6947 = _zz_6948;
  assign _zz_6948 = ($signed(_zz_6949) >>> _zz_775);
  assign _zz_6949 = _zz_6950;
  assign _zz_6950 = ($signed(data_mid_1_imag) - $signed(_zz_774));
  assign _zz_6951 = _zz_6952;
  assign _zz_6952 = ($signed(_zz_6953) >>> _zz_776);
  assign _zz_6953 = _zz_6954;
  assign _zz_6954 = ($signed(data_mid_1_real) + $signed(_zz_773));
  assign _zz_6955 = _zz_6956;
  assign _zz_6956 = ($signed(_zz_6957) >>> _zz_776);
  assign _zz_6957 = _zz_6958;
  assign _zz_6958 = ($signed(data_mid_1_imag) + $signed(_zz_774));
  assign _zz_6959 = ($signed(twiddle_factor_table_9_real) * $signed(data_mid_10_real));
  assign _zz_6960 = ($signed(twiddle_factor_table_9_imag) * $signed(data_mid_10_imag));
  assign _zz_6961 = fixTo_388_dout;
  assign _zz_6962 = ($signed(twiddle_factor_table_9_real) * $signed(data_mid_10_imag));
  assign _zz_6963 = ($signed(twiddle_factor_table_9_imag) * $signed(data_mid_10_real));
  assign _zz_6964 = fixTo_389_dout;
  assign _zz_6965 = _zz_6966;
  assign _zz_6966 = ($signed(_zz_6967) >>> _zz_779);
  assign _zz_6967 = _zz_6968;
  assign _zz_6968 = ($signed(data_mid_2_real) - $signed(_zz_777));
  assign _zz_6969 = _zz_6970;
  assign _zz_6970 = ($signed(_zz_6971) >>> _zz_779);
  assign _zz_6971 = _zz_6972;
  assign _zz_6972 = ($signed(data_mid_2_imag) - $signed(_zz_778));
  assign _zz_6973 = _zz_6974;
  assign _zz_6974 = ($signed(_zz_6975) >>> _zz_780);
  assign _zz_6975 = _zz_6976;
  assign _zz_6976 = ($signed(data_mid_2_real) + $signed(_zz_777));
  assign _zz_6977 = _zz_6978;
  assign _zz_6978 = ($signed(_zz_6979) >>> _zz_780);
  assign _zz_6979 = _zz_6980;
  assign _zz_6980 = ($signed(data_mid_2_imag) + $signed(_zz_778));
  assign _zz_6981 = ($signed(twiddle_factor_table_10_real) * $signed(data_mid_11_real));
  assign _zz_6982 = ($signed(twiddle_factor_table_10_imag) * $signed(data_mid_11_imag));
  assign _zz_6983 = fixTo_390_dout;
  assign _zz_6984 = ($signed(twiddle_factor_table_10_real) * $signed(data_mid_11_imag));
  assign _zz_6985 = ($signed(twiddle_factor_table_10_imag) * $signed(data_mid_11_real));
  assign _zz_6986 = fixTo_391_dout;
  assign _zz_6987 = _zz_6988;
  assign _zz_6988 = ($signed(_zz_6989) >>> _zz_783);
  assign _zz_6989 = _zz_6990;
  assign _zz_6990 = ($signed(data_mid_3_real) - $signed(_zz_781));
  assign _zz_6991 = _zz_6992;
  assign _zz_6992 = ($signed(_zz_6993) >>> _zz_783);
  assign _zz_6993 = _zz_6994;
  assign _zz_6994 = ($signed(data_mid_3_imag) - $signed(_zz_782));
  assign _zz_6995 = _zz_6996;
  assign _zz_6996 = ($signed(_zz_6997) >>> _zz_784);
  assign _zz_6997 = _zz_6998;
  assign _zz_6998 = ($signed(data_mid_3_real) + $signed(_zz_781));
  assign _zz_6999 = _zz_7000;
  assign _zz_7000 = ($signed(_zz_7001) >>> _zz_784);
  assign _zz_7001 = _zz_7002;
  assign _zz_7002 = ($signed(data_mid_3_imag) + $signed(_zz_782));
  assign _zz_7003 = ($signed(twiddle_factor_table_11_real) * $signed(data_mid_12_real));
  assign _zz_7004 = ($signed(twiddle_factor_table_11_imag) * $signed(data_mid_12_imag));
  assign _zz_7005 = fixTo_392_dout;
  assign _zz_7006 = ($signed(twiddle_factor_table_11_real) * $signed(data_mid_12_imag));
  assign _zz_7007 = ($signed(twiddle_factor_table_11_imag) * $signed(data_mid_12_real));
  assign _zz_7008 = fixTo_393_dout;
  assign _zz_7009 = _zz_7010;
  assign _zz_7010 = ($signed(_zz_7011) >>> _zz_787);
  assign _zz_7011 = _zz_7012;
  assign _zz_7012 = ($signed(data_mid_4_real) - $signed(_zz_785));
  assign _zz_7013 = _zz_7014;
  assign _zz_7014 = ($signed(_zz_7015) >>> _zz_787);
  assign _zz_7015 = _zz_7016;
  assign _zz_7016 = ($signed(data_mid_4_imag) - $signed(_zz_786));
  assign _zz_7017 = _zz_7018;
  assign _zz_7018 = ($signed(_zz_7019) >>> _zz_788);
  assign _zz_7019 = _zz_7020;
  assign _zz_7020 = ($signed(data_mid_4_real) + $signed(_zz_785));
  assign _zz_7021 = _zz_7022;
  assign _zz_7022 = ($signed(_zz_7023) >>> _zz_788);
  assign _zz_7023 = _zz_7024;
  assign _zz_7024 = ($signed(data_mid_4_imag) + $signed(_zz_786));
  assign _zz_7025 = ($signed(twiddle_factor_table_12_real) * $signed(data_mid_13_real));
  assign _zz_7026 = ($signed(twiddle_factor_table_12_imag) * $signed(data_mid_13_imag));
  assign _zz_7027 = fixTo_394_dout;
  assign _zz_7028 = ($signed(twiddle_factor_table_12_real) * $signed(data_mid_13_imag));
  assign _zz_7029 = ($signed(twiddle_factor_table_12_imag) * $signed(data_mid_13_real));
  assign _zz_7030 = fixTo_395_dout;
  assign _zz_7031 = _zz_7032;
  assign _zz_7032 = ($signed(_zz_7033) >>> _zz_791);
  assign _zz_7033 = _zz_7034;
  assign _zz_7034 = ($signed(data_mid_5_real) - $signed(_zz_789));
  assign _zz_7035 = _zz_7036;
  assign _zz_7036 = ($signed(_zz_7037) >>> _zz_791);
  assign _zz_7037 = _zz_7038;
  assign _zz_7038 = ($signed(data_mid_5_imag) - $signed(_zz_790));
  assign _zz_7039 = _zz_7040;
  assign _zz_7040 = ($signed(_zz_7041) >>> _zz_792);
  assign _zz_7041 = _zz_7042;
  assign _zz_7042 = ($signed(data_mid_5_real) + $signed(_zz_789));
  assign _zz_7043 = _zz_7044;
  assign _zz_7044 = ($signed(_zz_7045) >>> _zz_792);
  assign _zz_7045 = _zz_7046;
  assign _zz_7046 = ($signed(data_mid_5_imag) + $signed(_zz_790));
  assign _zz_7047 = ($signed(twiddle_factor_table_13_real) * $signed(data_mid_14_real));
  assign _zz_7048 = ($signed(twiddle_factor_table_13_imag) * $signed(data_mid_14_imag));
  assign _zz_7049 = fixTo_396_dout;
  assign _zz_7050 = ($signed(twiddle_factor_table_13_real) * $signed(data_mid_14_imag));
  assign _zz_7051 = ($signed(twiddle_factor_table_13_imag) * $signed(data_mid_14_real));
  assign _zz_7052 = fixTo_397_dout;
  assign _zz_7053 = _zz_7054;
  assign _zz_7054 = ($signed(_zz_7055) >>> _zz_795);
  assign _zz_7055 = _zz_7056;
  assign _zz_7056 = ($signed(data_mid_6_real) - $signed(_zz_793));
  assign _zz_7057 = _zz_7058;
  assign _zz_7058 = ($signed(_zz_7059) >>> _zz_795);
  assign _zz_7059 = _zz_7060;
  assign _zz_7060 = ($signed(data_mid_6_imag) - $signed(_zz_794));
  assign _zz_7061 = _zz_7062;
  assign _zz_7062 = ($signed(_zz_7063) >>> _zz_796);
  assign _zz_7063 = _zz_7064;
  assign _zz_7064 = ($signed(data_mid_6_real) + $signed(_zz_793));
  assign _zz_7065 = _zz_7066;
  assign _zz_7066 = ($signed(_zz_7067) >>> _zz_796);
  assign _zz_7067 = _zz_7068;
  assign _zz_7068 = ($signed(data_mid_6_imag) + $signed(_zz_794));
  assign _zz_7069 = ($signed(twiddle_factor_table_14_real) * $signed(data_mid_15_real));
  assign _zz_7070 = ($signed(twiddle_factor_table_14_imag) * $signed(data_mid_15_imag));
  assign _zz_7071 = fixTo_398_dout;
  assign _zz_7072 = ($signed(twiddle_factor_table_14_real) * $signed(data_mid_15_imag));
  assign _zz_7073 = ($signed(twiddle_factor_table_14_imag) * $signed(data_mid_15_real));
  assign _zz_7074 = fixTo_399_dout;
  assign _zz_7075 = _zz_7076;
  assign _zz_7076 = ($signed(_zz_7077) >>> _zz_799);
  assign _zz_7077 = _zz_7078;
  assign _zz_7078 = ($signed(data_mid_7_real) - $signed(_zz_797));
  assign _zz_7079 = _zz_7080;
  assign _zz_7080 = ($signed(_zz_7081) >>> _zz_799);
  assign _zz_7081 = _zz_7082;
  assign _zz_7082 = ($signed(data_mid_7_imag) - $signed(_zz_798));
  assign _zz_7083 = _zz_7084;
  assign _zz_7084 = ($signed(_zz_7085) >>> _zz_800);
  assign _zz_7085 = _zz_7086;
  assign _zz_7086 = ($signed(data_mid_7_real) + $signed(_zz_797));
  assign _zz_7087 = _zz_7088;
  assign _zz_7088 = ($signed(_zz_7089) >>> _zz_800);
  assign _zz_7089 = _zz_7090;
  assign _zz_7090 = ($signed(data_mid_7_imag) + $signed(_zz_798));
  assign _zz_7091 = ($signed(twiddle_factor_table_7_real) * $signed(data_mid_24_real));
  assign _zz_7092 = ($signed(twiddle_factor_table_7_imag) * $signed(data_mid_24_imag));
  assign _zz_7093 = fixTo_400_dout;
  assign _zz_7094 = ($signed(twiddle_factor_table_7_real) * $signed(data_mid_24_imag));
  assign _zz_7095 = ($signed(twiddle_factor_table_7_imag) * $signed(data_mid_24_real));
  assign _zz_7096 = fixTo_401_dout;
  assign _zz_7097 = _zz_7098;
  assign _zz_7098 = ($signed(_zz_7099) >>> _zz_803);
  assign _zz_7099 = _zz_7100;
  assign _zz_7100 = ($signed(data_mid_16_real) - $signed(_zz_801));
  assign _zz_7101 = _zz_7102;
  assign _zz_7102 = ($signed(_zz_7103) >>> _zz_803);
  assign _zz_7103 = _zz_7104;
  assign _zz_7104 = ($signed(data_mid_16_imag) - $signed(_zz_802));
  assign _zz_7105 = _zz_7106;
  assign _zz_7106 = ($signed(_zz_7107) >>> _zz_804);
  assign _zz_7107 = _zz_7108;
  assign _zz_7108 = ($signed(data_mid_16_real) + $signed(_zz_801));
  assign _zz_7109 = _zz_7110;
  assign _zz_7110 = ($signed(_zz_7111) >>> _zz_804);
  assign _zz_7111 = _zz_7112;
  assign _zz_7112 = ($signed(data_mid_16_imag) + $signed(_zz_802));
  assign _zz_7113 = ($signed(twiddle_factor_table_8_real) * $signed(data_mid_25_real));
  assign _zz_7114 = ($signed(twiddle_factor_table_8_imag) * $signed(data_mid_25_imag));
  assign _zz_7115 = fixTo_402_dout;
  assign _zz_7116 = ($signed(twiddle_factor_table_8_real) * $signed(data_mid_25_imag));
  assign _zz_7117 = ($signed(twiddle_factor_table_8_imag) * $signed(data_mid_25_real));
  assign _zz_7118 = fixTo_403_dout;
  assign _zz_7119 = _zz_7120;
  assign _zz_7120 = ($signed(_zz_7121) >>> _zz_807);
  assign _zz_7121 = _zz_7122;
  assign _zz_7122 = ($signed(data_mid_17_real) - $signed(_zz_805));
  assign _zz_7123 = _zz_7124;
  assign _zz_7124 = ($signed(_zz_7125) >>> _zz_807);
  assign _zz_7125 = _zz_7126;
  assign _zz_7126 = ($signed(data_mid_17_imag) - $signed(_zz_806));
  assign _zz_7127 = _zz_7128;
  assign _zz_7128 = ($signed(_zz_7129) >>> _zz_808);
  assign _zz_7129 = _zz_7130;
  assign _zz_7130 = ($signed(data_mid_17_real) + $signed(_zz_805));
  assign _zz_7131 = _zz_7132;
  assign _zz_7132 = ($signed(_zz_7133) >>> _zz_808);
  assign _zz_7133 = _zz_7134;
  assign _zz_7134 = ($signed(data_mid_17_imag) + $signed(_zz_806));
  assign _zz_7135 = ($signed(twiddle_factor_table_9_real) * $signed(data_mid_26_real));
  assign _zz_7136 = ($signed(twiddle_factor_table_9_imag) * $signed(data_mid_26_imag));
  assign _zz_7137 = fixTo_404_dout;
  assign _zz_7138 = ($signed(twiddle_factor_table_9_real) * $signed(data_mid_26_imag));
  assign _zz_7139 = ($signed(twiddle_factor_table_9_imag) * $signed(data_mid_26_real));
  assign _zz_7140 = fixTo_405_dout;
  assign _zz_7141 = _zz_7142;
  assign _zz_7142 = ($signed(_zz_7143) >>> _zz_811);
  assign _zz_7143 = _zz_7144;
  assign _zz_7144 = ($signed(data_mid_18_real) - $signed(_zz_809));
  assign _zz_7145 = _zz_7146;
  assign _zz_7146 = ($signed(_zz_7147) >>> _zz_811);
  assign _zz_7147 = _zz_7148;
  assign _zz_7148 = ($signed(data_mid_18_imag) - $signed(_zz_810));
  assign _zz_7149 = _zz_7150;
  assign _zz_7150 = ($signed(_zz_7151) >>> _zz_812);
  assign _zz_7151 = _zz_7152;
  assign _zz_7152 = ($signed(data_mid_18_real) + $signed(_zz_809));
  assign _zz_7153 = _zz_7154;
  assign _zz_7154 = ($signed(_zz_7155) >>> _zz_812);
  assign _zz_7155 = _zz_7156;
  assign _zz_7156 = ($signed(data_mid_18_imag) + $signed(_zz_810));
  assign _zz_7157 = ($signed(twiddle_factor_table_10_real) * $signed(data_mid_27_real));
  assign _zz_7158 = ($signed(twiddle_factor_table_10_imag) * $signed(data_mid_27_imag));
  assign _zz_7159 = fixTo_406_dout;
  assign _zz_7160 = ($signed(twiddle_factor_table_10_real) * $signed(data_mid_27_imag));
  assign _zz_7161 = ($signed(twiddle_factor_table_10_imag) * $signed(data_mid_27_real));
  assign _zz_7162 = fixTo_407_dout;
  assign _zz_7163 = _zz_7164;
  assign _zz_7164 = ($signed(_zz_7165) >>> _zz_815);
  assign _zz_7165 = _zz_7166;
  assign _zz_7166 = ($signed(data_mid_19_real) - $signed(_zz_813));
  assign _zz_7167 = _zz_7168;
  assign _zz_7168 = ($signed(_zz_7169) >>> _zz_815);
  assign _zz_7169 = _zz_7170;
  assign _zz_7170 = ($signed(data_mid_19_imag) - $signed(_zz_814));
  assign _zz_7171 = _zz_7172;
  assign _zz_7172 = ($signed(_zz_7173) >>> _zz_816);
  assign _zz_7173 = _zz_7174;
  assign _zz_7174 = ($signed(data_mid_19_real) + $signed(_zz_813));
  assign _zz_7175 = _zz_7176;
  assign _zz_7176 = ($signed(_zz_7177) >>> _zz_816);
  assign _zz_7177 = _zz_7178;
  assign _zz_7178 = ($signed(data_mid_19_imag) + $signed(_zz_814));
  assign _zz_7179 = ($signed(twiddle_factor_table_11_real) * $signed(data_mid_28_real));
  assign _zz_7180 = ($signed(twiddle_factor_table_11_imag) * $signed(data_mid_28_imag));
  assign _zz_7181 = fixTo_408_dout;
  assign _zz_7182 = ($signed(twiddle_factor_table_11_real) * $signed(data_mid_28_imag));
  assign _zz_7183 = ($signed(twiddle_factor_table_11_imag) * $signed(data_mid_28_real));
  assign _zz_7184 = fixTo_409_dout;
  assign _zz_7185 = _zz_7186;
  assign _zz_7186 = ($signed(_zz_7187) >>> _zz_819);
  assign _zz_7187 = _zz_7188;
  assign _zz_7188 = ($signed(data_mid_20_real) - $signed(_zz_817));
  assign _zz_7189 = _zz_7190;
  assign _zz_7190 = ($signed(_zz_7191) >>> _zz_819);
  assign _zz_7191 = _zz_7192;
  assign _zz_7192 = ($signed(data_mid_20_imag) - $signed(_zz_818));
  assign _zz_7193 = _zz_7194;
  assign _zz_7194 = ($signed(_zz_7195) >>> _zz_820);
  assign _zz_7195 = _zz_7196;
  assign _zz_7196 = ($signed(data_mid_20_real) + $signed(_zz_817));
  assign _zz_7197 = _zz_7198;
  assign _zz_7198 = ($signed(_zz_7199) >>> _zz_820);
  assign _zz_7199 = _zz_7200;
  assign _zz_7200 = ($signed(data_mid_20_imag) + $signed(_zz_818));
  assign _zz_7201 = ($signed(twiddle_factor_table_12_real) * $signed(data_mid_29_real));
  assign _zz_7202 = ($signed(twiddle_factor_table_12_imag) * $signed(data_mid_29_imag));
  assign _zz_7203 = fixTo_410_dout;
  assign _zz_7204 = ($signed(twiddle_factor_table_12_real) * $signed(data_mid_29_imag));
  assign _zz_7205 = ($signed(twiddle_factor_table_12_imag) * $signed(data_mid_29_real));
  assign _zz_7206 = fixTo_411_dout;
  assign _zz_7207 = _zz_7208;
  assign _zz_7208 = ($signed(_zz_7209) >>> _zz_823);
  assign _zz_7209 = _zz_7210;
  assign _zz_7210 = ($signed(data_mid_21_real) - $signed(_zz_821));
  assign _zz_7211 = _zz_7212;
  assign _zz_7212 = ($signed(_zz_7213) >>> _zz_823);
  assign _zz_7213 = _zz_7214;
  assign _zz_7214 = ($signed(data_mid_21_imag) - $signed(_zz_822));
  assign _zz_7215 = _zz_7216;
  assign _zz_7216 = ($signed(_zz_7217) >>> _zz_824);
  assign _zz_7217 = _zz_7218;
  assign _zz_7218 = ($signed(data_mid_21_real) + $signed(_zz_821));
  assign _zz_7219 = _zz_7220;
  assign _zz_7220 = ($signed(_zz_7221) >>> _zz_824);
  assign _zz_7221 = _zz_7222;
  assign _zz_7222 = ($signed(data_mid_21_imag) + $signed(_zz_822));
  assign _zz_7223 = ($signed(twiddle_factor_table_13_real) * $signed(data_mid_30_real));
  assign _zz_7224 = ($signed(twiddle_factor_table_13_imag) * $signed(data_mid_30_imag));
  assign _zz_7225 = fixTo_412_dout;
  assign _zz_7226 = ($signed(twiddle_factor_table_13_real) * $signed(data_mid_30_imag));
  assign _zz_7227 = ($signed(twiddle_factor_table_13_imag) * $signed(data_mid_30_real));
  assign _zz_7228 = fixTo_413_dout;
  assign _zz_7229 = _zz_7230;
  assign _zz_7230 = ($signed(_zz_7231) >>> _zz_827);
  assign _zz_7231 = _zz_7232;
  assign _zz_7232 = ($signed(data_mid_22_real) - $signed(_zz_825));
  assign _zz_7233 = _zz_7234;
  assign _zz_7234 = ($signed(_zz_7235) >>> _zz_827);
  assign _zz_7235 = _zz_7236;
  assign _zz_7236 = ($signed(data_mid_22_imag) - $signed(_zz_826));
  assign _zz_7237 = _zz_7238;
  assign _zz_7238 = ($signed(_zz_7239) >>> _zz_828);
  assign _zz_7239 = _zz_7240;
  assign _zz_7240 = ($signed(data_mid_22_real) + $signed(_zz_825));
  assign _zz_7241 = _zz_7242;
  assign _zz_7242 = ($signed(_zz_7243) >>> _zz_828);
  assign _zz_7243 = _zz_7244;
  assign _zz_7244 = ($signed(data_mid_22_imag) + $signed(_zz_826));
  assign _zz_7245 = ($signed(twiddle_factor_table_14_real) * $signed(data_mid_31_real));
  assign _zz_7246 = ($signed(twiddle_factor_table_14_imag) * $signed(data_mid_31_imag));
  assign _zz_7247 = fixTo_414_dout;
  assign _zz_7248 = ($signed(twiddle_factor_table_14_real) * $signed(data_mid_31_imag));
  assign _zz_7249 = ($signed(twiddle_factor_table_14_imag) * $signed(data_mid_31_real));
  assign _zz_7250 = fixTo_415_dout;
  assign _zz_7251 = _zz_7252;
  assign _zz_7252 = ($signed(_zz_7253) >>> _zz_831);
  assign _zz_7253 = _zz_7254;
  assign _zz_7254 = ($signed(data_mid_23_real) - $signed(_zz_829));
  assign _zz_7255 = _zz_7256;
  assign _zz_7256 = ($signed(_zz_7257) >>> _zz_831);
  assign _zz_7257 = _zz_7258;
  assign _zz_7258 = ($signed(data_mid_23_imag) - $signed(_zz_830));
  assign _zz_7259 = _zz_7260;
  assign _zz_7260 = ($signed(_zz_7261) >>> _zz_832);
  assign _zz_7261 = _zz_7262;
  assign _zz_7262 = ($signed(data_mid_23_real) + $signed(_zz_829));
  assign _zz_7263 = _zz_7264;
  assign _zz_7264 = ($signed(_zz_7265) >>> _zz_832);
  assign _zz_7265 = _zz_7266;
  assign _zz_7266 = ($signed(data_mid_23_imag) + $signed(_zz_830));
  assign _zz_7267 = ($signed(twiddle_factor_table_7_real) * $signed(data_mid_40_real));
  assign _zz_7268 = ($signed(twiddle_factor_table_7_imag) * $signed(data_mid_40_imag));
  assign _zz_7269 = fixTo_416_dout;
  assign _zz_7270 = ($signed(twiddle_factor_table_7_real) * $signed(data_mid_40_imag));
  assign _zz_7271 = ($signed(twiddle_factor_table_7_imag) * $signed(data_mid_40_real));
  assign _zz_7272 = fixTo_417_dout;
  assign _zz_7273 = _zz_7274;
  assign _zz_7274 = ($signed(_zz_7275) >>> _zz_835);
  assign _zz_7275 = _zz_7276;
  assign _zz_7276 = ($signed(data_mid_32_real) - $signed(_zz_833));
  assign _zz_7277 = _zz_7278;
  assign _zz_7278 = ($signed(_zz_7279) >>> _zz_835);
  assign _zz_7279 = _zz_7280;
  assign _zz_7280 = ($signed(data_mid_32_imag) - $signed(_zz_834));
  assign _zz_7281 = _zz_7282;
  assign _zz_7282 = ($signed(_zz_7283) >>> _zz_836);
  assign _zz_7283 = _zz_7284;
  assign _zz_7284 = ($signed(data_mid_32_real) + $signed(_zz_833));
  assign _zz_7285 = _zz_7286;
  assign _zz_7286 = ($signed(_zz_7287) >>> _zz_836);
  assign _zz_7287 = _zz_7288;
  assign _zz_7288 = ($signed(data_mid_32_imag) + $signed(_zz_834));
  assign _zz_7289 = ($signed(twiddle_factor_table_8_real) * $signed(data_mid_41_real));
  assign _zz_7290 = ($signed(twiddle_factor_table_8_imag) * $signed(data_mid_41_imag));
  assign _zz_7291 = fixTo_418_dout;
  assign _zz_7292 = ($signed(twiddle_factor_table_8_real) * $signed(data_mid_41_imag));
  assign _zz_7293 = ($signed(twiddle_factor_table_8_imag) * $signed(data_mid_41_real));
  assign _zz_7294 = fixTo_419_dout;
  assign _zz_7295 = _zz_7296;
  assign _zz_7296 = ($signed(_zz_7297) >>> _zz_839);
  assign _zz_7297 = _zz_7298;
  assign _zz_7298 = ($signed(data_mid_33_real) - $signed(_zz_837));
  assign _zz_7299 = _zz_7300;
  assign _zz_7300 = ($signed(_zz_7301) >>> _zz_839);
  assign _zz_7301 = _zz_7302;
  assign _zz_7302 = ($signed(data_mid_33_imag) - $signed(_zz_838));
  assign _zz_7303 = _zz_7304;
  assign _zz_7304 = ($signed(_zz_7305) >>> _zz_840);
  assign _zz_7305 = _zz_7306;
  assign _zz_7306 = ($signed(data_mid_33_real) + $signed(_zz_837));
  assign _zz_7307 = _zz_7308;
  assign _zz_7308 = ($signed(_zz_7309) >>> _zz_840);
  assign _zz_7309 = _zz_7310;
  assign _zz_7310 = ($signed(data_mid_33_imag) + $signed(_zz_838));
  assign _zz_7311 = ($signed(twiddle_factor_table_9_real) * $signed(data_mid_42_real));
  assign _zz_7312 = ($signed(twiddle_factor_table_9_imag) * $signed(data_mid_42_imag));
  assign _zz_7313 = fixTo_420_dout;
  assign _zz_7314 = ($signed(twiddle_factor_table_9_real) * $signed(data_mid_42_imag));
  assign _zz_7315 = ($signed(twiddle_factor_table_9_imag) * $signed(data_mid_42_real));
  assign _zz_7316 = fixTo_421_dout;
  assign _zz_7317 = _zz_7318;
  assign _zz_7318 = ($signed(_zz_7319) >>> _zz_843);
  assign _zz_7319 = _zz_7320;
  assign _zz_7320 = ($signed(data_mid_34_real) - $signed(_zz_841));
  assign _zz_7321 = _zz_7322;
  assign _zz_7322 = ($signed(_zz_7323) >>> _zz_843);
  assign _zz_7323 = _zz_7324;
  assign _zz_7324 = ($signed(data_mid_34_imag) - $signed(_zz_842));
  assign _zz_7325 = _zz_7326;
  assign _zz_7326 = ($signed(_zz_7327) >>> _zz_844);
  assign _zz_7327 = _zz_7328;
  assign _zz_7328 = ($signed(data_mid_34_real) + $signed(_zz_841));
  assign _zz_7329 = _zz_7330;
  assign _zz_7330 = ($signed(_zz_7331) >>> _zz_844);
  assign _zz_7331 = _zz_7332;
  assign _zz_7332 = ($signed(data_mid_34_imag) + $signed(_zz_842));
  assign _zz_7333 = ($signed(twiddle_factor_table_10_real) * $signed(data_mid_43_real));
  assign _zz_7334 = ($signed(twiddle_factor_table_10_imag) * $signed(data_mid_43_imag));
  assign _zz_7335 = fixTo_422_dout;
  assign _zz_7336 = ($signed(twiddle_factor_table_10_real) * $signed(data_mid_43_imag));
  assign _zz_7337 = ($signed(twiddle_factor_table_10_imag) * $signed(data_mid_43_real));
  assign _zz_7338 = fixTo_423_dout;
  assign _zz_7339 = _zz_7340;
  assign _zz_7340 = ($signed(_zz_7341) >>> _zz_847);
  assign _zz_7341 = _zz_7342;
  assign _zz_7342 = ($signed(data_mid_35_real) - $signed(_zz_845));
  assign _zz_7343 = _zz_7344;
  assign _zz_7344 = ($signed(_zz_7345) >>> _zz_847);
  assign _zz_7345 = _zz_7346;
  assign _zz_7346 = ($signed(data_mid_35_imag) - $signed(_zz_846));
  assign _zz_7347 = _zz_7348;
  assign _zz_7348 = ($signed(_zz_7349) >>> _zz_848);
  assign _zz_7349 = _zz_7350;
  assign _zz_7350 = ($signed(data_mid_35_real) + $signed(_zz_845));
  assign _zz_7351 = _zz_7352;
  assign _zz_7352 = ($signed(_zz_7353) >>> _zz_848);
  assign _zz_7353 = _zz_7354;
  assign _zz_7354 = ($signed(data_mid_35_imag) + $signed(_zz_846));
  assign _zz_7355 = ($signed(twiddle_factor_table_11_real) * $signed(data_mid_44_real));
  assign _zz_7356 = ($signed(twiddle_factor_table_11_imag) * $signed(data_mid_44_imag));
  assign _zz_7357 = fixTo_424_dout;
  assign _zz_7358 = ($signed(twiddle_factor_table_11_real) * $signed(data_mid_44_imag));
  assign _zz_7359 = ($signed(twiddle_factor_table_11_imag) * $signed(data_mid_44_real));
  assign _zz_7360 = fixTo_425_dout;
  assign _zz_7361 = _zz_7362;
  assign _zz_7362 = ($signed(_zz_7363) >>> _zz_851);
  assign _zz_7363 = _zz_7364;
  assign _zz_7364 = ($signed(data_mid_36_real) - $signed(_zz_849));
  assign _zz_7365 = _zz_7366;
  assign _zz_7366 = ($signed(_zz_7367) >>> _zz_851);
  assign _zz_7367 = _zz_7368;
  assign _zz_7368 = ($signed(data_mid_36_imag) - $signed(_zz_850));
  assign _zz_7369 = _zz_7370;
  assign _zz_7370 = ($signed(_zz_7371) >>> _zz_852);
  assign _zz_7371 = _zz_7372;
  assign _zz_7372 = ($signed(data_mid_36_real) + $signed(_zz_849));
  assign _zz_7373 = _zz_7374;
  assign _zz_7374 = ($signed(_zz_7375) >>> _zz_852);
  assign _zz_7375 = _zz_7376;
  assign _zz_7376 = ($signed(data_mid_36_imag) + $signed(_zz_850));
  assign _zz_7377 = ($signed(twiddle_factor_table_12_real) * $signed(data_mid_45_real));
  assign _zz_7378 = ($signed(twiddle_factor_table_12_imag) * $signed(data_mid_45_imag));
  assign _zz_7379 = fixTo_426_dout;
  assign _zz_7380 = ($signed(twiddle_factor_table_12_real) * $signed(data_mid_45_imag));
  assign _zz_7381 = ($signed(twiddle_factor_table_12_imag) * $signed(data_mid_45_real));
  assign _zz_7382 = fixTo_427_dout;
  assign _zz_7383 = _zz_7384;
  assign _zz_7384 = ($signed(_zz_7385) >>> _zz_855);
  assign _zz_7385 = _zz_7386;
  assign _zz_7386 = ($signed(data_mid_37_real) - $signed(_zz_853));
  assign _zz_7387 = _zz_7388;
  assign _zz_7388 = ($signed(_zz_7389) >>> _zz_855);
  assign _zz_7389 = _zz_7390;
  assign _zz_7390 = ($signed(data_mid_37_imag) - $signed(_zz_854));
  assign _zz_7391 = _zz_7392;
  assign _zz_7392 = ($signed(_zz_7393) >>> _zz_856);
  assign _zz_7393 = _zz_7394;
  assign _zz_7394 = ($signed(data_mid_37_real) + $signed(_zz_853));
  assign _zz_7395 = _zz_7396;
  assign _zz_7396 = ($signed(_zz_7397) >>> _zz_856);
  assign _zz_7397 = _zz_7398;
  assign _zz_7398 = ($signed(data_mid_37_imag) + $signed(_zz_854));
  assign _zz_7399 = ($signed(twiddle_factor_table_13_real) * $signed(data_mid_46_real));
  assign _zz_7400 = ($signed(twiddle_factor_table_13_imag) * $signed(data_mid_46_imag));
  assign _zz_7401 = fixTo_428_dout;
  assign _zz_7402 = ($signed(twiddle_factor_table_13_real) * $signed(data_mid_46_imag));
  assign _zz_7403 = ($signed(twiddle_factor_table_13_imag) * $signed(data_mid_46_real));
  assign _zz_7404 = fixTo_429_dout;
  assign _zz_7405 = _zz_7406;
  assign _zz_7406 = ($signed(_zz_7407) >>> _zz_859);
  assign _zz_7407 = _zz_7408;
  assign _zz_7408 = ($signed(data_mid_38_real) - $signed(_zz_857));
  assign _zz_7409 = _zz_7410;
  assign _zz_7410 = ($signed(_zz_7411) >>> _zz_859);
  assign _zz_7411 = _zz_7412;
  assign _zz_7412 = ($signed(data_mid_38_imag) - $signed(_zz_858));
  assign _zz_7413 = _zz_7414;
  assign _zz_7414 = ($signed(_zz_7415) >>> _zz_860);
  assign _zz_7415 = _zz_7416;
  assign _zz_7416 = ($signed(data_mid_38_real) + $signed(_zz_857));
  assign _zz_7417 = _zz_7418;
  assign _zz_7418 = ($signed(_zz_7419) >>> _zz_860);
  assign _zz_7419 = _zz_7420;
  assign _zz_7420 = ($signed(data_mid_38_imag) + $signed(_zz_858));
  assign _zz_7421 = ($signed(twiddle_factor_table_14_real) * $signed(data_mid_47_real));
  assign _zz_7422 = ($signed(twiddle_factor_table_14_imag) * $signed(data_mid_47_imag));
  assign _zz_7423 = fixTo_430_dout;
  assign _zz_7424 = ($signed(twiddle_factor_table_14_real) * $signed(data_mid_47_imag));
  assign _zz_7425 = ($signed(twiddle_factor_table_14_imag) * $signed(data_mid_47_real));
  assign _zz_7426 = fixTo_431_dout;
  assign _zz_7427 = _zz_7428;
  assign _zz_7428 = ($signed(_zz_7429) >>> _zz_863);
  assign _zz_7429 = _zz_7430;
  assign _zz_7430 = ($signed(data_mid_39_real) - $signed(_zz_861));
  assign _zz_7431 = _zz_7432;
  assign _zz_7432 = ($signed(_zz_7433) >>> _zz_863);
  assign _zz_7433 = _zz_7434;
  assign _zz_7434 = ($signed(data_mid_39_imag) - $signed(_zz_862));
  assign _zz_7435 = _zz_7436;
  assign _zz_7436 = ($signed(_zz_7437) >>> _zz_864);
  assign _zz_7437 = _zz_7438;
  assign _zz_7438 = ($signed(data_mid_39_real) + $signed(_zz_861));
  assign _zz_7439 = _zz_7440;
  assign _zz_7440 = ($signed(_zz_7441) >>> _zz_864);
  assign _zz_7441 = _zz_7442;
  assign _zz_7442 = ($signed(data_mid_39_imag) + $signed(_zz_862));
  assign _zz_7443 = ($signed(twiddle_factor_table_7_real) * $signed(data_mid_56_real));
  assign _zz_7444 = ($signed(twiddle_factor_table_7_imag) * $signed(data_mid_56_imag));
  assign _zz_7445 = fixTo_432_dout;
  assign _zz_7446 = ($signed(twiddle_factor_table_7_real) * $signed(data_mid_56_imag));
  assign _zz_7447 = ($signed(twiddle_factor_table_7_imag) * $signed(data_mid_56_real));
  assign _zz_7448 = fixTo_433_dout;
  assign _zz_7449 = _zz_7450;
  assign _zz_7450 = ($signed(_zz_7451) >>> _zz_867);
  assign _zz_7451 = _zz_7452;
  assign _zz_7452 = ($signed(data_mid_48_real) - $signed(_zz_865));
  assign _zz_7453 = _zz_7454;
  assign _zz_7454 = ($signed(_zz_7455) >>> _zz_867);
  assign _zz_7455 = _zz_7456;
  assign _zz_7456 = ($signed(data_mid_48_imag) - $signed(_zz_866));
  assign _zz_7457 = _zz_7458;
  assign _zz_7458 = ($signed(_zz_7459) >>> _zz_868);
  assign _zz_7459 = _zz_7460;
  assign _zz_7460 = ($signed(data_mid_48_real) + $signed(_zz_865));
  assign _zz_7461 = _zz_7462;
  assign _zz_7462 = ($signed(_zz_7463) >>> _zz_868);
  assign _zz_7463 = _zz_7464;
  assign _zz_7464 = ($signed(data_mid_48_imag) + $signed(_zz_866));
  assign _zz_7465 = ($signed(twiddle_factor_table_8_real) * $signed(data_mid_57_real));
  assign _zz_7466 = ($signed(twiddle_factor_table_8_imag) * $signed(data_mid_57_imag));
  assign _zz_7467 = fixTo_434_dout;
  assign _zz_7468 = ($signed(twiddle_factor_table_8_real) * $signed(data_mid_57_imag));
  assign _zz_7469 = ($signed(twiddle_factor_table_8_imag) * $signed(data_mid_57_real));
  assign _zz_7470 = fixTo_435_dout;
  assign _zz_7471 = _zz_7472;
  assign _zz_7472 = ($signed(_zz_7473) >>> _zz_871);
  assign _zz_7473 = _zz_7474;
  assign _zz_7474 = ($signed(data_mid_49_real) - $signed(_zz_869));
  assign _zz_7475 = _zz_7476;
  assign _zz_7476 = ($signed(_zz_7477) >>> _zz_871);
  assign _zz_7477 = _zz_7478;
  assign _zz_7478 = ($signed(data_mid_49_imag) - $signed(_zz_870));
  assign _zz_7479 = _zz_7480;
  assign _zz_7480 = ($signed(_zz_7481) >>> _zz_872);
  assign _zz_7481 = _zz_7482;
  assign _zz_7482 = ($signed(data_mid_49_real) + $signed(_zz_869));
  assign _zz_7483 = _zz_7484;
  assign _zz_7484 = ($signed(_zz_7485) >>> _zz_872);
  assign _zz_7485 = _zz_7486;
  assign _zz_7486 = ($signed(data_mid_49_imag) + $signed(_zz_870));
  assign _zz_7487 = ($signed(twiddle_factor_table_9_real) * $signed(data_mid_58_real));
  assign _zz_7488 = ($signed(twiddle_factor_table_9_imag) * $signed(data_mid_58_imag));
  assign _zz_7489 = fixTo_436_dout;
  assign _zz_7490 = ($signed(twiddle_factor_table_9_real) * $signed(data_mid_58_imag));
  assign _zz_7491 = ($signed(twiddle_factor_table_9_imag) * $signed(data_mid_58_real));
  assign _zz_7492 = fixTo_437_dout;
  assign _zz_7493 = _zz_7494;
  assign _zz_7494 = ($signed(_zz_7495) >>> _zz_875);
  assign _zz_7495 = _zz_7496;
  assign _zz_7496 = ($signed(data_mid_50_real) - $signed(_zz_873));
  assign _zz_7497 = _zz_7498;
  assign _zz_7498 = ($signed(_zz_7499) >>> _zz_875);
  assign _zz_7499 = _zz_7500;
  assign _zz_7500 = ($signed(data_mid_50_imag) - $signed(_zz_874));
  assign _zz_7501 = _zz_7502;
  assign _zz_7502 = ($signed(_zz_7503) >>> _zz_876);
  assign _zz_7503 = _zz_7504;
  assign _zz_7504 = ($signed(data_mid_50_real) + $signed(_zz_873));
  assign _zz_7505 = _zz_7506;
  assign _zz_7506 = ($signed(_zz_7507) >>> _zz_876);
  assign _zz_7507 = _zz_7508;
  assign _zz_7508 = ($signed(data_mid_50_imag) + $signed(_zz_874));
  assign _zz_7509 = ($signed(twiddle_factor_table_10_real) * $signed(data_mid_59_real));
  assign _zz_7510 = ($signed(twiddle_factor_table_10_imag) * $signed(data_mid_59_imag));
  assign _zz_7511 = fixTo_438_dout;
  assign _zz_7512 = ($signed(twiddle_factor_table_10_real) * $signed(data_mid_59_imag));
  assign _zz_7513 = ($signed(twiddle_factor_table_10_imag) * $signed(data_mid_59_real));
  assign _zz_7514 = fixTo_439_dout;
  assign _zz_7515 = _zz_7516;
  assign _zz_7516 = ($signed(_zz_7517) >>> _zz_879);
  assign _zz_7517 = _zz_7518;
  assign _zz_7518 = ($signed(data_mid_51_real) - $signed(_zz_877));
  assign _zz_7519 = _zz_7520;
  assign _zz_7520 = ($signed(_zz_7521) >>> _zz_879);
  assign _zz_7521 = _zz_7522;
  assign _zz_7522 = ($signed(data_mid_51_imag) - $signed(_zz_878));
  assign _zz_7523 = _zz_7524;
  assign _zz_7524 = ($signed(_zz_7525) >>> _zz_880);
  assign _zz_7525 = _zz_7526;
  assign _zz_7526 = ($signed(data_mid_51_real) + $signed(_zz_877));
  assign _zz_7527 = _zz_7528;
  assign _zz_7528 = ($signed(_zz_7529) >>> _zz_880);
  assign _zz_7529 = _zz_7530;
  assign _zz_7530 = ($signed(data_mid_51_imag) + $signed(_zz_878));
  assign _zz_7531 = ($signed(twiddle_factor_table_11_real) * $signed(data_mid_60_real));
  assign _zz_7532 = ($signed(twiddle_factor_table_11_imag) * $signed(data_mid_60_imag));
  assign _zz_7533 = fixTo_440_dout;
  assign _zz_7534 = ($signed(twiddle_factor_table_11_real) * $signed(data_mid_60_imag));
  assign _zz_7535 = ($signed(twiddle_factor_table_11_imag) * $signed(data_mid_60_real));
  assign _zz_7536 = fixTo_441_dout;
  assign _zz_7537 = _zz_7538;
  assign _zz_7538 = ($signed(_zz_7539) >>> _zz_883);
  assign _zz_7539 = _zz_7540;
  assign _zz_7540 = ($signed(data_mid_52_real) - $signed(_zz_881));
  assign _zz_7541 = _zz_7542;
  assign _zz_7542 = ($signed(_zz_7543) >>> _zz_883);
  assign _zz_7543 = _zz_7544;
  assign _zz_7544 = ($signed(data_mid_52_imag) - $signed(_zz_882));
  assign _zz_7545 = _zz_7546;
  assign _zz_7546 = ($signed(_zz_7547) >>> _zz_884);
  assign _zz_7547 = _zz_7548;
  assign _zz_7548 = ($signed(data_mid_52_real) + $signed(_zz_881));
  assign _zz_7549 = _zz_7550;
  assign _zz_7550 = ($signed(_zz_7551) >>> _zz_884);
  assign _zz_7551 = _zz_7552;
  assign _zz_7552 = ($signed(data_mid_52_imag) + $signed(_zz_882));
  assign _zz_7553 = ($signed(twiddle_factor_table_12_real) * $signed(data_mid_61_real));
  assign _zz_7554 = ($signed(twiddle_factor_table_12_imag) * $signed(data_mid_61_imag));
  assign _zz_7555 = fixTo_442_dout;
  assign _zz_7556 = ($signed(twiddle_factor_table_12_real) * $signed(data_mid_61_imag));
  assign _zz_7557 = ($signed(twiddle_factor_table_12_imag) * $signed(data_mid_61_real));
  assign _zz_7558 = fixTo_443_dout;
  assign _zz_7559 = _zz_7560;
  assign _zz_7560 = ($signed(_zz_7561) >>> _zz_887);
  assign _zz_7561 = _zz_7562;
  assign _zz_7562 = ($signed(data_mid_53_real) - $signed(_zz_885));
  assign _zz_7563 = _zz_7564;
  assign _zz_7564 = ($signed(_zz_7565) >>> _zz_887);
  assign _zz_7565 = _zz_7566;
  assign _zz_7566 = ($signed(data_mid_53_imag) - $signed(_zz_886));
  assign _zz_7567 = _zz_7568;
  assign _zz_7568 = ($signed(_zz_7569) >>> _zz_888);
  assign _zz_7569 = _zz_7570;
  assign _zz_7570 = ($signed(data_mid_53_real) + $signed(_zz_885));
  assign _zz_7571 = _zz_7572;
  assign _zz_7572 = ($signed(_zz_7573) >>> _zz_888);
  assign _zz_7573 = _zz_7574;
  assign _zz_7574 = ($signed(data_mid_53_imag) + $signed(_zz_886));
  assign _zz_7575 = ($signed(twiddle_factor_table_13_real) * $signed(data_mid_62_real));
  assign _zz_7576 = ($signed(twiddle_factor_table_13_imag) * $signed(data_mid_62_imag));
  assign _zz_7577 = fixTo_444_dout;
  assign _zz_7578 = ($signed(twiddle_factor_table_13_real) * $signed(data_mid_62_imag));
  assign _zz_7579 = ($signed(twiddle_factor_table_13_imag) * $signed(data_mid_62_real));
  assign _zz_7580 = fixTo_445_dout;
  assign _zz_7581 = _zz_7582;
  assign _zz_7582 = ($signed(_zz_7583) >>> _zz_891);
  assign _zz_7583 = _zz_7584;
  assign _zz_7584 = ($signed(data_mid_54_real) - $signed(_zz_889));
  assign _zz_7585 = _zz_7586;
  assign _zz_7586 = ($signed(_zz_7587) >>> _zz_891);
  assign _zz_7587 = _zz_7588;
  assign _zz_7588 = ($signed(data_mid_54_imag) - $signed(_zz_890));
  assign _zz_7589 = _zz_7590;
  assign _zz_7590 = ($signed(_zz_7591) >>> _zz_892);
  assign _zz_7591 = _zz_7592;
  assign _zz_7592 = ($signed(data_mid_54_real) + $signed(_zz_889));
  assign _zz_7593 = _zz_7594;
  assign _zz_7594 = ($signed(_zz_7595) >>> _zz_892);
  assign _zz_7595 = _zz_7596;
  assign _zz_7596 = ($signed(data_mid_54_imag) + $signed(_zz_890));
  assign _zz_7597 = ($signed(twiddle_factor_table_14_real) * $signed(data_mid_63_real));
  assign _zz_7598 = ($signed(twiddle_factor_table_14_imag) * $signed(data_mid_63_imag));
  assign _zz_7599 = fixTo_446_dout;
  assign _zz_7600 = ($signed(twiddle_factor_table_14_real) * $signed(data_mid_63_imag));
  assign _zz_7601 = ($signed(twiddle_factor_table_14_imag) * $signed(data_mid_63_real));
  assign _zz_7602 = fixTo_447_dout;
  assign _zz_7603 = _zz_7604;
  assign _zz_7604 = ($signed(_zz_7605) >>> _zz_895);
  assign _zz_7605 = _zz_7606;
  assign _zz_7606 = ($signed(data_mid_55_real) - $signed(_zz_893));
  assign _zz_7607 = _zz_7608;
  assign _zz_7608 = ($signed(_zz_7609) >>> _zz_895);
  assign _zz_7609 = _zz_7610;
  assign _zz_7610 = ($signed(data_mid_55_imag) - $signed(_zz_894));
  assign _zz_7611 = _zz_7612;
  assign _zz_7612 = ($signed(_zz_7613) >>> _zz_896);
  assign _zz_7613 = _zz_7614;
  assign _zz_7614 = ($signed(data_mid_55_real) + $signed(_zz_893));
  assign _zz_7615 = _zz_7616;
  assign _zz_7616 = ($signed(_zz_7617) >>> _zz_896);
  assign _zz_7617 = _zz_7618;
  assign _zz_7618 = ($signed(data_mid_55_imag) + $signed(_zz_894));
  assign _zz_7619 = ($signed(twiddle_factor_table_7_real) * $signed(data_mid_72_real));
  assign _zz_7620 = ($signed(twiddle_factor_table_7_imag) * $signed(data_mid_72_imag));
  assign _zz_7621 = fixTo_448_dout;
  assign _zz_7622 = ($signed(twiddle_factor_table_7_real) * $signed(data_mid_72_imag));
  assign _zz_7623 = ($signed(twiddle_factor_table_7_imag) * $signed(data_mid_72_real));
  assign _zz_7624 = fixTo_449_dout;
  assign _zz_7625 = _zz_7626;
  assign _zz_7626 = ($signed(_zz_7627) >>> _zz_899);
  assign _zz_7627 = _zz_7628;
  assign _zz_7628 = ($signed(data_mid_64_real) - $signed(_zz_897));
  assign _zz_7629 = _zz_7630;
  assign _zz_7630 = ($signed(_zz_7631) >>> _zz_899);
  assign _zz_7631 = _zz_7632;
  assign _zz_7632 = ($signed(data_mid_64_imag) - $signed(_zz_898));
  assign _zz_7633 = _zz_7634;
  assign _zz_7634 = ($signed(_zz_7635) >>> _zz_900);
  assign _zz_7635 = _zz_7636;
  assign _zz_7636 = ($signed(data_mid_64_real) + $signed(_zz_897));
  assign _zz_7637 = _zz_7638;
  assign _zz_7638 = ($signed(_zz_7639) >>> _zz_900);
  assign _zz_7639 = _zz_7640;
  assign _zz_7640 = ($signed(data_mid_64_imag) + $signed(_zz_898));
  assign _zz_7641 = ($signed(twiddle_factor_table_8_real) * $signed(data_mid_73_real));
  assign _zz_7642 = ($signed(twiddle_factor_table_8_imag) * $signed(data_mid_73_imag));
  assign _zz_7643 = fixTo_450_dout;
  assign _zz_7644 = ($signed(twiddle_factor_table_8_real) * $signed(data_mid_73_imag));
  assign _zz_7645 = ($signed(twiddle_factor_table_8_imag) * $signed(data_mid_73_real));
  assign _zz_7646 = fixTo_451_dout;
  assign _zz_7647 = _zz_7648;
  assign _zz_7648 = ($signed(_zz_7649) >>> _zz_903);
  assign _zz_7649 = _zz_7650;
  assign _zz_7650 = ($signed(data_mid_65_real) - $signed(_zz_901));
  assign _zz_7651 = _zz_7652;
  assign _zz_7652 = ($signed(_zz_7653) >>> _zz_903);
  assign _zz_7653 = _zz_7654;
  assign _zz_7654 = ($signed(data_mid_65_imag) - $signed(_zz_902));
  assign _zz_7655 = _zz_7656;
  assign _zz_7656 = ($signed(_zz_7657) >>> _zz_904);
  assign _zz_7657 = _zz_7658;
  assign _zz_7658 = ($signed(data_mid_65_real) + $signed(_zz_901));
  assign _zz_7659 = _zz_7660;
  assign _zz_7660 = ($signed(_zz_7661) >>> _zz_904);
  assign _zz_7661 = _zz_7662;
  assign _zz_7662 = ($signed(data_mid_65_imag) + $signed(_zz_902));
  assign _zz_7663 = ($signed(twiddle_factor_table_9_real) * $signed(data_mid_74_real));
  assign _zz_7664 = ($signed(twiddle_factor_table_9_imag) * $signed(data_mid_74_imag));
  assign _zz_7665 = fixTo_452_dout;
  assign _zz_7666 = ($signed(twiddle_factor_table_9_real) * $signed(data_mid_74_imag));
  assign _zz_7667 = ($signed(twiddle_factor_table_9_imag) * $signed(data_mid_74_real));
  assign _zz_7668 = fixTo_453_dout;
  assign _zz_7669 = _zz_7670;
  assign _zz_7670 = ($signed(_zz_7671) >>> _zz_907);
  assign _zz_7671 = _zz_7672;
  assign _zz_7672 = ($signed(data_mid_66_real) - $signed(_zz_905));
  assign _zz_7673 = _zz_7674;
  assign _zz_7674 = ($signed(_zz_7675) >>> _zz_907);
  assign _zz_7675 = _zz_7676;
  assign _zz_7676 = ($signed(data_mid_66_imag) - $signed(_zz_906));
  assign _zz_7677 = _zz_7678;
  assign _zz_7678 = ($signed(_zz_7679) >>> _zz_908);
  assign _zz_7679 = _zz_7680;
  assign _zz_7680 = ($signed(data_mid_66_real) + $signed(_zz_905));
  assign _zz_7681 = _zz_7682;
  assign _zz_7682 = ($signed(_zz_7683) >>> _zz_908);
  assign _zz_7683 = _zz_7684;
  assign _zz_7684 = ($signed(data_mid_66_imag) + $signed(_zz_906));
  assign _zz_7685 = ($signed(twiddle_factor_table_10_real) * $signed(data_mid_75_real));
  assign _zz_7686 = ($signed(twiddle_factor_table_10_imag) * $signed(data_mid_75_imag));
  assign _zz_7687 = fixTo_454_dout;
  assign _zz_7688 = ($signed(twiddle_factor_table_10_real) * $signed(data_mid_75_imag));
  assign _zz_7689 = ($signed(twiddle_factor_table_10_imag) * $signed(data_mid_75_real));
  assign _zz_7690 = fixTo_455_dout;
  assign _zz_7691 = _zz_7692;
  assign _zz_7692 = ($signed(_zz_7693) >>> _zz_911);
  assign _zz_7693 = _zz_7694;
  assign _zz_7694 = ($signed(data_mid_67_real) - $signed(_zz_909));
  assign _zz_7695 = _zz_7696;
  assign _zz_7696 = ($signed(_zz_7697) >>> _zz_911);
  assign _zz_7697 = _zz_7698;
  assign _zz_7698 = ($signed(data_mid_67_imag) - $signed(_zz_910));
  assign _zz_7699 = _zz_7700;
  assign _zz_7700 = ($signed(_zz_7701) >>> _zz_912);
  assign _zz_7701 = _zz_7702;
  assign _zz_7702 = ($signed(data_mid_67_real) + $signed(_zz_909));
  assign _zz_7703 = _zz_7704;
  assign _zz_7704 = ($signed(_zz_7705) >>> _zz_912);
  assign _zz_7705 = _zz_7706;
  assign _zz_7706 = ($signed(data_mid_67_imag) + $signed(_zz_910));
  assign _zz_7707 = ($signed(twiddle_factor_table_11_real) * $signed(data_mid_76_real));
  assign _zz_7708 = ($signed(twiddle_factor_table_11_imag) * $signed(data_mid_76_imag));
  assign _zz_7709 = fixTo_456_dout;
  assign _zz_7710 = ($signed(twiddle_factor_table_11_real) * $signed(data_mid_76_imag));
  assign _zz_7711 = ($signed(twiddle_factor_table_11_imag) * $signed(data_mid_76_real));
  assign _zz_7712 = fixTo_457_dout;
  assign _zz_7713 = _zz_7714;
  assign _zz_7714 = ($signed(_zz_7715) >>> _zz_915);
  assign _zz_7715 = _zz_7716;
  assign _zz_7716 = ($signed(data_mid_68_real) - $signed(_zz_913));
  assign _zz_7717 = _zz_7718;
  assign _zz_7718 = ($signed(_zz_7719) >>> _zz_915);
  assign _zz_7719 = _zz_7720;
  assign _zz_7720 = ($signed(data_mid_68_imag) - $signed(_zz_914));
  assign _zz_7721 = _zz_7722;
  assign _zz_7722 = ($signed(_zz_7723) >>> _zz_916);
  assign _zz_7723 = _zz_7724;
  assign _zz_7724 = ($signed(data_mid_68_real) + $signed(_zz_913));
  assign _zz_7725 = _zz_7726;
  assign _zz_7726 = ($signed(_zz_7727) >>> _zz_916);
  assign _zz_7727 = _zz_7728;
  assign _zz_7728 = ($signed(data_mid_68_imag) + $signed(_zz_914));
  assign _zz_7729 = ($signed(twiddle_factor_table_12_real) * $signed(data_mid_77_real));
  assign _zz_7730 = ($signed(twiddle_factor_table_12_imag) * $signed(data_mid_77_imag));
  assign _zz_7731 = fixTo_458_dout;
  assign _zz_7732 = ($signed(twiddle_factor_table_12_real) * $signed(data_mid_77_imag));
  assign _zz_7733 = ($signed(twiddle_factor_table_12_imag) * $signed(data_mid_77_real));
  assign _zz_7734 = fixTo_459_dout;
  assign _zz_7735 = _zz_7736;
  assign _zz_7736 = ($signed(_zz_7737) >>> _zz_919);
  assign _zz_7737 = _zz_7738;
  assign _zz_7738 = ($signed(data_mid_69_real) - $signed(_zz_917));
  assign _zz_7739 = _zz_7740;
  assign _zz_7740 = ($signed(_zz_7741) >>> _zz_919);
  assign _zz_7741 = _zz_7742;
  assign _zz_7742 = ($signed(data_mid_69_imag) - $signed(_zz_918));
  assign _zz_7743 = _zz_7744;
  assign _zz_7744 = ($signed(_zz_7745) >>> _zz_920);
  assign _zz_7745 = _zz_7746;
  assign _zz_7746 = ($signed(data_mid_69_real) + $signed(_zz_917));
  assign _zz_7747 = _zz_7748;
  assign _zz_7748 = ($signed(_zz_7749) >>> _zz_920);
  assign _zz_7749 = _zz_7750;
  assign _zz_7750 = ($signed(data_mid_69_imag) + $signed(_zz_918));
  assign _zz_7751 = ($signed(twiddle_factor_table_13_real) * $signed(data_mid_78_real));
  assign _zz_7752 = ($signed(twiddle_factor_table_13_imag) * $signed(data_mid_78_imag));
  assign _zz_7753 = fixTo_460_dout;
  assign _zz_7754 = ($signed(twiddle_factor_table_13_real) * $signed(data_mid_78_imag));
  assign _zz_7755 = ($signed(twiddle_factor_table_13_imag) * $signed(data_mid_78_real));
  assign _zz_7756 = fixTo_461_dout;
  assign _zz_7757 = _zz_7758;
  assign _zz_7758 = ($signed(_zz_7759) >>> _zz_923);
  assign _zz_7759 = _zz_7760;
  assign _zz_7760 = ($signed(data_mid_70_real) - $signed(_zz_921));
  assign _zz_7761 = _zz_7762;
  assign _zz_7762 = ($signed(_zz_7763) >>> _zz_923);
  assign _zz_7763 = _zz_7764;
  assign _zz_7764 = ($signed(data_mid_70_imag) - $signed(_zz_922));
  assign _zz_7765 = _zz_7766;
  assign _zz_7766 = ($signed(_zz_7767) >>> _zz_924);
  assign _zz_7767 = _zz_7768;
  assign _zz_7768 = ($signed(data_mid_70_real) + $signed(_zz_921));
  assign _zz_7769 = _zz_7770;
  assign _zz_7770 = ($signed(_zz_7771) >>> _zz_924);
  assign _zz_7771 = _zz_7772;
  assign _zz_7772 = ($signed(data_mid_70_imag) + $signed(_zz_922));
  assign _zz_7773 = ($signed(twiddle_factor_table_14_real) * $signed(data_mid_79_real));
  assign _zz_7774 = ($signed(twiddle_factor_table_14_imag) * $signed(data_mid_79_imag));
  assign _zz_7775 = fixTo_462_dout;
  assign _zz_7776 = ($signed(twiddle_factor_table_14_real) * $signed(data_mid_79_imag));
  assign _zz_7777 = ($signed(twiddle_factor_table_14_imag) * $signed(data_mid_79_real));
  assign _zz_7778 = fixTo_463_dout;
  assign _zz_7779 = _zz_7780;
  assign _zz_7780 = ($signed(_zz_7781) >>> _zz_927);
  assign _zz_7781 = _zz_7782;
  assign _zz_7782 = ($signed(data_mid_71_real) - $signed(_zz_925));
  assign _zz_7783 = _zz_7784;
  assign _zz_7784 = ($signed(_zz_7785) >>> _zz_927);
  assign _zz_7785 = _zz_7786;
  assign _zz_7786 = ($signed(data_mid_71_imag) - $signed(_zz_926));
  assign _zz_7787 = _zz_7788;
  assign _zz_7788 = ($signed(_zz_7789) >>> _zz_928);
  assign _zz_7789 = _zz_7790;
  assign _zz_7790 = ($signed(data_mid_71_real) + $signed(_zz_925));
  assign _zz_7791 = _zz_7792;
  assign _zz_7792 = ($signed(_zz_7793) >>> _zz_928);
  assign _zz_7793 = _zz_7794;
  assign _zz_7794 = ($signed(data_mid_71_imag) + $signed(_zz_926));
  assign _zz_7795 = ($signed(twiddle_factor_table_7_real) * $signed(data_mid_88_real));
  assign _zz_7796 = ($signed(twiddle_factor_table_7_imag) * $signed(data_mid_88_imag));
  assign _zz_7797 = fixTo_464_dout;
  assign _zz_7798 = ($signed(twiddle_factor_table_7_real) * $signed(data_mid_88_imag));
  assign _zz_7799 = ($signed(twiddle_factor_table_7_imag) * $signed(data_mid_88_real));
  assign _zz_7800 = fixTo_465_dout;
  assign _zz_7801 = _zz_7802;
  assign _zz_7802 = ($signed(_zz_7803) >>> _zz_931);
  assign _zz_7803 = _zz_7804;
  assign _zz_7804 = ($signed(data_mid_80_real) - $signed(_zz_929));
  assign _zz_7805 = _zz_7806;
  assign _zz_7806 = ($signed(_zz_7807) >>> _zz_931);
  assign _zz_7807 = _zz_7808;
  assign _zz_7808 = ($signed(data_mid_80_imag) - $signed(_zz_930));
  assign _zz_7809 = _zz_7810;
  assign _zz_7810 = ($signed(_zz_7811) >>> _zz_932);
  assign _zz_7811 = _zz_7812;
  assign _zz_7812 = ($signed(data_mid_80_real) + $signed(_zz_929));
  assign _zz_7813 = _zz_7814;
  assign _zz_7814 = ($signed(_zz_7815) >>> _zz_932);
  assign _zz_7815 = _zz_7816;
  assign _zz_7816 = ($signed(data_mid_80_imag) + $signed(_zz_930));
  assign _zz_7817 = ($signed(twiddle_factor_table_8_real) * $signed(data_mid_89_real));
  assign _zz_7818 = ($signed(twiddle_factor_table_8_imag) * $signed(data_mid_89_imag));
  assign _zz_7819 = fixTo_466_dout;
  assign _zz_7820 = ($signed(twiddle_factor_table_8_real) * $signed(data_mid_89_imag));
  assign _zz_7821 = ($signed(twiddle_factor_table_8_imag) * $signed(data_mid_89_real));
  assign _zz_7822 = fixTo_467_dout;
  assign _zz_7823 = _zz_7824;
  assign _zz_7824 = ($signed(_zz_7825) >>> _zz_935);
  assign _zz_7825 = _zz_7826;
  assign _zz_7826 = ($signed(data_mid_81_real) - $signed(_zz_933));
  assign _zz_7827 = _zz_7828;
  assign _zz_7828 = ($signed(_zz_7829) >>> _zz_935);
  assign _zz_7829 = _zz_7830;
  assign _zz_7830 = ($signed(data_mid_81_imag) - $signed(_zz_934));
  assign _zz_7831 = _zz_7832;
  assign _zz_7832 = ($signed(_zz_7833) >>> _zz_936);
  assign _zz_7833 = _zz_7834;
  assign _zz_7834 = ($signed(data_mid_81_real) + $signed(_zz_933));
  assign _zz_7835 = _zz_7836;
  assign _zz_7836 = ($signed(_zz_7837) >>> _zz_936);
  assign _zz_7837 = _zz_7838;
  assign _zz_7838 = ($signed(data_mid_81_imag) + $signed(_zz_934));
  assign _zz_7839 = ($signed(twiddle_factor_table_9_real) * $signed(data_mid_90_real));
  assign _zz_7840 = ($signed(twiddle_factor_table_9_imag) * $signed(data_mid_90_imag));
  assign _zz_7841 = fixTo_468_dout;
  assign _zz_7842 = ($signed(twiddle_factor_table_9_real) * $signed(data_mid_90_imag));
  assign _zz_7843 = ($signed(twiddle_factor_table_9_imag) * $signed(data_mid_90_real));
  assign _zz_7844 = fixTo_469_dout;
  assign _zz_7845 = _zz_7846;
  assign _zz_7846 = ($signed(_zz_7847) >>> _zz_939);
  assign _zz_7847 = _zz_7848;
  assign _zz_7848 = ($signed(data_mid_82_real) - $signed(_zz_937));
  assign _zz_7849 = _zz_7850;
  assign _zz_7850 = ($signed(_zz_7851) >>> _zz_939);
  assign _zz_7851 = _zz_7852;
  assign _zz_7852 = ($signed(data_mid_82_imag) - $signed(_zz_938));
  assign _zz_7853 = _zz_7854;
  assign _zz_7854 = ($signed(_zz_7855) >>> _zz_940);
  assign _zz_7855 = _zz_7856;
  assign _zz_7856 = ($signed(data_mid_82_real) + $signed(_zz_937));
  assign _zz_7857 = _zz_7858;
  assign _zz_7858 = ($signed(_zz_7859) >>> _zz_940);
  assign _zz_7859 = _zz_7860;
  assign _zz_7860 = ($signed(data_mid_82_imag) + $signed(_zz_938));
  assign _zz_7861 = ($signed(twiddle_factor_table_10_real) * $signed(data_mid_91_real));
  assign _zz_7862 = ($signed(twiddle_factor_table_10_imag) * $signed(data_mid_91_imag));
  assign _zz_7863 = fixTo_470_dout;
  assign _zz_7864 = ($signed(twiddle_factor_table_10_real) * $signed(data_mid_91_imag));
  assign _zz_7865 = ($signed(twiddle_factor_table_10_imag) * $signed(data_mid_91_real));
  assign _zz_7866 = fixTo_471_dout;
  assign _zz_7867 = _zz_7868;
  assign _zz_7868 = ($signed(_zz_7869) >>> _zz_943);
  assign _zz_7869 = _zz_7870;
  assign _zz_7870 = ($signed(data_mid_83_real) - $signed(_zz_941));
  assign _zz_7871 = _zz_7872;
  assign _zz_7872 = ($signed(_zz_7873) >>> _zz_943);
  assign _zz_7873 = _zz_7874;
  assign _zz_7874 = ($signed(data_mid_83_imag) - $signed(_zz_942));
  assign _zz_7875 = _zz_7876;
  assign _zz_7876 = ($signed(_zz_7877) >>> _zz_944);
  assign _zz_7877 = _zz_7878;
  assign _zz_7878 = ($signed(data_mid_83_real) + $signed(_zz_941));
  assign _zz_7879 = _zz_7880;
  assign _zz_7880 = ($signed(_zz_7881) >>> _zz_944);
  assign _zz_7881 = _zz_7882;
  assign _zz_7882 = ($signed(data_mid_83_imag) + $signed(_zz_942));
  assign _zz_7883 = ($signed(twiddle_factor_table_11_real) * $signed(data_mid_92_real));
  assign _zz_7884 = ($signed(twiddle_factor_table_11_imag) * $signed(data_mid_92_imag));
  assign _zz_7885 = fixTo_472_dout;
  assign _zz_7886 = ($signed(twiddle_factor_table_11_real) * $signed(data_mid_92_imag));
  assign _zz_7887 = ($signed(twiddle_factor_table_11_imag) * $signed(data_mid_92_real));
  assign _zz_7888 = fixTo_473_dout;
  assign _zz_7889 = _zz_7890;
  assign _zz_7890 = ($signed(_zz_7891) >>> _zz_947);
  assign _zz_7891 = _zz_7892;
  assign _zz_7892 = ($signed(data_mid_84_real) - $signed(_zz_945));
  assign _zz_7893 = _zz_7894;
  assign _zz_7894 = ($signed(_zz_7895) >>> _zz_947);
  assign _zz_7895 = _zz_7896;
  assign _zz_7896 = ($signed(data_mid_84_imag) - $signed(_zz_946));
  assign _zz_7897 = _zz_7898;
  assign _zz_7898 = ($signed(_zz_7899) >>> _zz_948);
  assign _zz_7899 = _zz_7900;
  assign _zz_7900 = ($signed(data_mid_84_real) + $signed(_zz_945));
  assign _zz_7901 = _zz_7902;
  assign _zz_7902 = ($signed(_zz_7903) >>> _zz_948);
  assign _zz_7903 = _zz_7904;
  assign _zz_7904 = ($signed(data_mid_84_imag) + $signed(_zz_946));
  assign _zz_7905 = ($signed(twiddle_factor_table_12_real) * $signed(data_mid_93_real));
  assign _zz_7906 = ($signed(twiddle_factor_table_12_imag) * $signed(data_mid_93_imag));
  assign _zz_7907 = fixTo_474_dout;
  assign _zz_7908 = ($signed(twiddle_factor_table_12_real) * $signed(data_mid_93_imag));
  assign _zz_7909 = ($signed(twiddle_factor_table_12_imag) * $signed(data_mid_93_real));
  assign _zz_7910 = fixTo_475_dout;
  assign _zz_7911 = _zz_7912;
  assign _zz_7912 = ($signed(_zz_7913) >>> _zz_951);
  assign _zz_7913 = _zz_7914;
  assign _zz_7914 = ($signed(data_mid_85_real) - $signed(_zz_949));
  assign _zz_7915 = _zz_7916;
  assign _zz_7916 = ($signed(_zz_7917) >>> _zz_951);
  assign _zz_7917 = _zz_7918;
  assign _zz_7918 = ($signed(data_mid_85_imag) - $signed(_zz_950));
  assign _zz_7919 = _zz_7920;
  assign _zz_7920 = ($signed(_zz_7921) >>> _zz_952);
  assign _zz_7921 = _zz_7922;
  assign _zz_7922 = ($signed(data_mid_85_real) + $signed(_zz_949));
  assign _zz_7923 = _zz_7924;
  assign _zz_7924 = ($signed(_zz_7925) >>> _zz_952);
  assign _zz_7925 = _zz_7926;
  assign _zz_7926 = ($signed(data_mid_85_imag) + $signed(_zz_950));
  assign _zz_7927 = ($signed(twiddle_factor_table_13_real) * $signed(data_mid_94_real));
  assign _zz_7928 = ($signed(twiddle_factor_table_13_imag) * $signed(data_mid_94_imag));
  assign _zz_7929 = fixTo_476_dout;
  assign _zz_7930 = ($signed(twiddle_factor_table_13_real) * $signed(data_mid_94_imag));
  assign _zz_7931 = ($signed(twiddle_factor_table_13_imag) * $signed(data_mid_94_real));
  assign _zz_7932 = fixTo_477_dout;
  assign _zz_7933 = _zz_7934;
  assign _zz_7934 = ($signed(_zz_7935) >>> _zz_955);
  assign _zz_7935 = _zz_7936;
  assign _zz_7936 = ($signed(data_mid_86_real) - $signed(_zz_953));
  assign _zz_7937 = _zz_7938;
  assign _zz_7938 = ($signed(_zz_7939) >>> _zz_955);
  assign _zz_7939 = _zz_7940;
  assign _zz_7940 = ($signed(data_mid_86_imag) - $signed(_zz_954));
  assign _zz_7941 = _zz_7942;
  assign _zz_7942 = ($signed(_zz_7943) >>> _zz_956);
  assign _zz_7943 = _zz_7944;
  assign _zz_7944 = ($signed(data_mid_86_real) + $signed(_zz_953));
  assign _zz_7945 = _zz_7946;
  assign _zz_7946 = ($signed(_zz_7947) >>> _zz_956);
  assign _zz_7947 = _zz_7948;
  assign _zz_7948 = ($signed(data_mid_86_imag) + $signed(_zz_954));
  assign _zz_7949 = ($signed(twiddle_factor_table_14_real) * $signed(data_mid_95_real));
  assign _zz_7950 = ($signed(twiddle_factor_table_14_imag) * $signed(data_mid_95_imag));
  assign _zz_7951 = fixTo_478_dout;
  assign _zz_7952 = ($signed(twiddle_factor_table_14_real) * $signed(data_mid_95_imag));
  assign _zz_7953 = ($signed(twiddle_factor_table_14_imag) * $signed(data_mid_95_real));
  assign _zz_7954 = fixTo_479_dout;
  assign _zz_7955 = _zz_7956;
  assign _zz_7956 = ($signed(_zz_7957) >>> _zz_959);
  assign _zz_7957 = _zz_7958;
  assign _zz_7958 = ($signed(data_mid_87_real) - $signed(_zz_957));
  assign _zz_7959 = _zz_7960;
  assign _zz_7960 = ($signed(_zz_7961) >>> _zz_959);
  assign _zz_7961 = _zz_7962;
  assign _zz_7962 = ($signed(data_mid_87_imag) - $signed(_zz_958));
  assign _zz_7963 = _zz_7964;
  assign _zz_7964 = ($signed(_zz_7965) >>> _zz_960);
  assign _zz_7965 = _zz_7966;
  assign _zz_7966 = ($signed(data_mid_87_real) + $signed(_zz_957));
  assign _zz_7967 = _zz_7968;
  assign _zz_7968 = ($signed(_zz_7969) >>> _zz_960);
  assign _zz_7969 = _zz_7970;
  assign _zz_7970 = ($signed(data_mid_87_imag) + $signed(_zz_958));
  assign _zz_7971 = ($signed(twiddle_factor_table_7_real) * $signed(data_mid_104_real));
  assign _zz_7972 = ($signed(twiddle_factor_table_7_imag) * $signed(data_mid_104_imag));
  assign _zz_7973 = fixTo_480_dout;
  assign _zz_7974 = ($signed(twiddle_factor_table_7_real) * $signed(data_mid_104_imag));
  assign _zz_7975 = ($signed(twiddle_factor_table_7_imag) * $signed(data_mid_104_real));
  assign _zz_7976 = fixTo_481_dout;
  assign _zz_7977 = _zz_7978;
  assign _zz_7978 = ($signed(_zz_7979) >>> _zz_963);
  assign _zz_7979 = _zz_7980;
  assign _zz_7980 = ($signed(data_mid_96_real) - $signed(_zz_961));
  assign _zz_7981 = _zz_7982;
  assign _zz_7982 = ($signed(_zz_7983) >>> _zz_963);
  assign _zz_7983 = _zz_7984;
  assign _zz_7984 = ($signed(data_mid_96_imag) - $signed(_zz_962));
  assign _zz_7985 = _zz_7986;
  assign _zz_7986 = ($signed(_zz_7987) >>> _zz_964);
  assign _zz_7987 = _zz_7988;
  assign _zz_7988 = ($signed(data_mid_96_real) + $signed(_zz_961));
  assign _zz_7989 = _zz_7990;
  assign _zz_7990 = ($signed(_zz_7991) >>> _zz_964);
  assign _zz_7991 = _zz_7992;
  assign _zz_7992 = ($signed(data_mid_96_imag) + $signed(_zz_962));
  assign _zz_7993 = ($signed(twiddle_factor_table_8_real) * $signed(data_mid_105_real));
  assign _zz_7994 = ($signed(twiddle_factor_table_8_imag) * $signed(data_mid_105_imag));
  assign _zz_7995 = fixTo_482_dout;
  assign _zz_7996 = ($signed(twiddle_factor_table_8_real) * $signed(data_mid_105_imag));
  assign _zz_7997 = ($signed(twiddle_factor_table_8_imag) * $signed(data_mid_105_real));
  assign _zz_7998 = fixTo_483_dout;
  assign _zz_7999 = _zz_8000;
  assign _zz_8000 = ($signed(_zz_8001) >>> _zz_967);
  assign _zz_8001 = _zz_8002;
  assign _zz_8002 = ($signed(data_mid_97_real) - $signed(_zz_965));
  assign _zz_8003 = _zz_8004;
  assign _zz_8004 = ($signed(_zz_8005) >>> _zz_967);
  assign _zz_8005 = _zz_8006;
  assign _zz_8006 = ($signed(data_mid_97_imag) - $signed(_zz_966));
  assign _zz_8007 = _zz_8008;
  assign _zz_8008 = ($signed(_zz_8009) >>> _zz_968);
  assign _zz_8009 = _zz_8010;
  assign _zz_8010 = ($signed(data_mid_97_real) + $signed(_zz_965));
  assign _zz_8011 = _zz_8012;
  assign _zz_8012 = ($signed(_zz_8013) >>> _zz_968);
  assign _zz_8013 = _zz_8014;
  assign _zz_8014 = ($signed(data_mid_97_imag) + $signed(_zz_966));
  assign _zz_8015 = ($signed(twiddle_factor_table_9_real) * $signed(data_mid_106_real));
  assign _zz_8016 = ($signed(twiddle_factor_table_9_imag) * $signed(data_mid_106_imag));
  assign _zz_8017 = fixTo_484_dout;
  assign _zz_8018 = ($signed(twiddle_factor_table_9_real) * $signed(data_mid_106_imag));
  assign _zz_8019 = ($signed(twiddle_factor_table_9_imag) * $signed(data_mid_106_real));
  assign _zz_8020 = fixTo_485_dout;
  assign _zz_8021 = _zz_8022;
  assign _zz_8022 = ($signed(_zz_8023) >>> _zz_971);
  assign _zz_8023 = _zz_8024;
  assign _zz_8024 = ($signed(data_mid_98_real) - $signed(_zz_969));
  assign _zz_8025 = _zz_8026;
  assign _zz_8026 = ($signed(_zz_8027) >>> _zz_971);
  assign _zz_8027 = _zz_8028;
  assign _zz_8028 = ($signed(data_mid_98_imag) - $signed(_zz_970));
  assign _zz_8029 = _zz_8030;
  assign _zz_8030 = ($signed(_zz_8031) >>> _zz_972);
  assign _zz_8031 = _zz_8032;
  assign _zz_8032 = ($signed(data_mid_98_real) + $signed(_zz_969));
  assign _zz_8033 = _zz_8034;
  assign _zz_8034 = ($signed(_zz_8035) >>> _zz_972);
  assign _zz_8035 = _zz_8036;
  assign _zz_8036 = ($signed(data_mid_98_imag) + $signed(_zz_970));
  assign _zz_8037 = ($signed(twiddle_factor_table_10_real) * $signed(data_mid_107_real));
  assign _zz_8038 = ($signed(twiddle_factor_table_10_imag) * $signed(data_mid_107_imag));
  assign _zz_8039 = fixTo_486_dout;
  assign _zz_8040 = ($signed(twiddle_factor_table_10_real) * $signed(data_mid_107_imag));
  assign _zz_8041 = ($signed(twiddle_factor_table_10_imag) * $signed(data_mid_107_real));
  assign _zz_8042 = fixTo_487_dout;
  assign _zz_8043 = _zz_8044;
  assign _zz_8044 = ($signed(_zz_8045) >>> _zz_975);
  assign _zz_8045 = _zz_8046;
  assign _zz_8046 = ($signed(data_mid_99_real) - $signed(_zz_973));
  assign _zz_8047 = _zz_8048;
  assign _zz_8048 = ($signed(_zz_8049) >>> _zz_975);
  assign _zz_8049 = _zz_8050;
  assign _zz_8050 = ($signed(data_mid_99_imag) - $signed(_zz_974));
  assign _zz_8051 = _zz_8052;
  assign _zz_8052 = ($signed(_zz_8053) >>> _zz_976);
  assign _zz_8053 = _zz_8054;
  assign _zz_8054 = ($signed(data_mid_99_real) + $signed(_zz_973));
  assign _zz_8055 = _zz_8056;
  assign _zz_8056 = ($signed(_zz_8057) >>> _zz_976);
  assign _zz_8057 = _zz_8058;
  assign _zz_8058 = ($signed(data_mid_99_imag) + $signed(_zz_974));
  assign _zz_8059 = ($signed(twiddle_factor_table_11_real) * $signed(data_mid_108_real));
  assign _zz_8060 = ($signed(twiddle_factor_table_11_imag) * $signed(data_mid_108_imag));
  assign _zz_8061 = fixTo_488_dout;
  assign _zz_8062 = ($signed(twiddle_factor_table_11_real) * $signed(data_mid_108_imag));
  assign _zz_8063 = ($signed(twiddle_factor_table_11_imag) * $signed(data_mid_108_real));
  assign _zz_8064 = fixTo_489_dout;
  assign _zz_8065 = _zz_8066;
  assign _zz_8066 = ($signed(_zz_8067) >>> _zz_979);
  assign _zz_8067 = _zz_8068;
  assign _zz_8068 = ($signed(data_mid_100_real) - $signed(_zz_977));
  assign _zz_8069 = _zz_8070;
  assign _zz_8070 = ($signed(_zz_8071) >>> _zz_979);
  assign _zz_8071 = _zz_8072;
  assign _zz_8072 = ($signed(data_mid_100_imag) - $signed(_zz_978));
  assign _zz_8073 = _zz_8074;
  assign _zz_8074 = ($signed(_zz_8075) >>> _zz_980);
  assign _zz_8075 = _zz_8076;
  assign _zz_8076 = ($signed(data_mid_100_real) + $signed(_zz_977));
  assign _zz_8077 = _zz_8078;
  assign _zz_8078 = ($signed(_zz_8079) >>> _zz_980);
  assign _zz_8079 = _zz_8080;
  assign _zz_8080 = ($signed(data_mid_100_imag) + $signed(_zz_978));
  assign _zz_8081 = ($signed(twiddle_factor_table_12_real) * $signed(data_mid_109_real));
  assign _zz_8082 = ($signed(twiddle_factor_table_12_imag) * $signed(data_mid_109_imag));
  assign _zz_8083 = fixTo_490_dout;
  assign _zz_8084 = ($signed(twiddle_factor_table_12_real) * $signed(data_mid_109_imag));
  assign _zz_8085 = ($signed(twiddle_factor_table_12_imag) * $signed(data_mid_109_real));
  assign _zz_8086 = fixTo_491_dout;
  assign _zz_8087 = _zz_8088;
  assign _zz_8088 = ($signed(_zz_8089) >>> _zz_983);
  assign _zz_8089 = _zz_8090;
  assign _zz_8090 = ($signed(data_mid_101_real) - $signed(_zz_981));
  assign _zz_8091 = _zz_8092;
  assign _zz_8092 = ($signed(_zz_8093) >>> _zz_983);
  assign _zz_8093 = _zz_8094;
  assign _zz_8094 = ($signed(data_mid_101_imag) - $signed(_zz_982));
  assign _zz_8095 = _zz_8096;
  assign _zz_8096 = ($signed(_zz_8097) >>> _zz_984);
  assign _zz_8097 = _zz_8098;
  assign _zz_8098 = ($signed(data_mid_101_real) + $signed(_zz_981));
  assign _zz_8099 = _zz_8100;
  assign _zz_8100 = ($signed(_zz_8101) >>> _zz_984);
  assign _zz_8101 = _zz_8102;
  assign _zz_8102 = ($signed(data_mid_101_imag) + $signed(_zz_982));
  assign _zz_8103 = ($signed(twiddle_factor_table_13_real) * $signed(data_mid_110_real));
  assign _zz_8104 = ($signed(twiddle_factor_table_13_imag) * $signed(data_mid_110_imag));
  assign _zz_8105 = fixTo_492_dout;
  assign _zz_8106 = ($signed(twiddle_factor_table_13_real) * $signed(data_mid_110_imag));
  assign _zz_8107 = ($signed(twiddle_factor_table_13_imag) * $signed(data_mid_110_real));
  assign _zz_8108 = fixTo_493_dout;
  assign _zz_8109 = _zz_8110;
  assign _zz_8110 = ($signed(_zz_8111) >>> _zz_987);
  assign _zz_8111 = _zz_8112;
  assign _zz_8112 = ($signed(data_mid_102_real) - $signed(_zz_985));
  assign _zz_8113 = _zz_8114;
  assign _zz_8114 = ($signed(_zz_8115) >>> _zz_987);
  assign _zz_8115 = _zz_8116;
  assign _zz_8116 = ($signed(data_mid_102_imag) - $signed(_zz_986));
  assign _zz_8117 = _zz_8118;
  assign _zz_8118 = ($signed(_zz_8119) >>> _zz_988);
  assign _zz_8119 = _zz_8120;
  assign _zz_8120 = ($signed(data_mid_102_real) + $signed(_zz_985));
  assign _zz_8121 = _zz_8122;
  assign _zz_8122 = ($signed(_zz_8123) >>> _zz_988);
  assign _zz_8123 = _zz_8124;
  assign _zz_8124 = ($signed(data_mid_102_imag) + $signed(_zz_986));
  assign _zz_8125 = ($signed(twiddle_factor_table_14_real) * $signed(data_mid_111_real));
  assign _zz_8126 = ($signed(twiddle_factor_table_14_imag) * $signed(data_mid_111_imag));
  assign _zz_8127 = fixTo_494_dout;
  assign _zz_8128 = ($signed(twiddle_factor_table_14_real) * $signed(data_mid_111_imag));
  assign _zz_8129 = ($signed(twiddle_factor_table_14_imag) * $signed(data_mid_111_real));
  assign _zz_8130 = fixTo_495_dout;
  assign _zz_8131 = _zz_8132;
  assign _zz_8132 = ($signed(_zz_8133) >>> _zz_991);
  assign _zz_8133 = _zz_8134;
  assign _zz_8134 = ($signed(data_mid_103_real) - $signed(_zz_989));
  assign _zz_8135 = _zz_8136;
  assign _zz_8136 = ($signed(_zz_8137) >>> _zz_991);
  assign _zz_8137 = _zz_8138;
  assign _zz_8138 = ($signed(data_mid_103_imag) - $signed(_zz_990));
  assign _zz_8139 = _zz_8140;
  assign _zz_8140 = ($signed(_zz_8141) >>> _zz_992);
  assign _zz_8141 = _zz_8142;
  assign _zz_8142 = ($signed(data_mid_103_real) + $signed(_zz_989));
  assign _zz_8143 = _zz_8144;
  assign _zz_8144 = ($signed(_zz_8145) >>> _zz_992);
  assign _zz_8145 = _zz_8146;
  assign _zz_8146 = ($signed(data_mid_103_imag) + $signed(_zz_990));
  assign _zz_8147 = ($signed(twiddle_factor_table_7_real) * $signed(data_mid_120_real));
  assign _zz_8148 = ($signed(twiddle_factor_table_7_imag) * $signed(data_mid_120_imag));
  assign _zz_8149 = fixTo_496_dout;
  assign _zz_8150 = ($signed(twiddle_factor_table_7_real) * $signed(data_mid_120_imag));
  assign _zz_8151 = ($signed(twiddle_factor_table_7_imag) * $signed(data_mid_120_real));
  assign _zz_8152 = fixTo_497_dout;
  assign _zz_8153 = _zz_8154;
  assign _zz_8154 = ($signed(_zz_8155) >>> _zz_995);
  assign _zz_8155 = _zz_8156;
  assign _zz_8156 = ($signed(data_mid_112_real) - $signed(_zz_993));
  assign _zz_8157 = _zz_8158;
  assign _zz_8158 = ($signed(_zz_8159) >>> _zz_995);
  assign _zz_8159 = _zz_8160;
  assign _zz_8160 = ($signed(data_mid_112_imag) - $signed(_zz_994));
  assign _zz_8161 = _zz_8162;
  assign _zz_8162 = ($signed(_zz_8163) >>> _zz_996);
  assign _zz_8163 = _zz_8164;
  assign _zz_8164 = ($signed(data_mid_112_real) + $signed(_zz_993));
  assign _zz_8165 = _zz_8166;
  assign _zz_8166 = ($signed(_zz_8167) >>> _zz_996);
  assign _zz_8167 = _zz_8168;
  assign _zz_8168 = ($signed(data_mid_112_imag) + $signed(_zz_994));
  assign _zz_8169 = ($signed(twiddle_factor_table_8_real) * $signed(data_mid_121_real));
  assign _zz_8170 = ($signed(twiddle_factor_table_8_imag) * $signed(data_mid_121_imag));
  assign _zz_8171 = fixTo_498_dout;
  assign _zz_8172 = ($signed(twiddle_factor_table_8_real) * $signed(data_mid_121_imag));
  assign _zz_8173 = ($signed(twiddle_factor_table_8_imag) * $signed(data_mid_121_real));
  assign _zz_8174 = fixTo_499_dout;
  assign _zz_8175 = _zz_8176;
  assign _zz_8176 = ($signed(_zz_8177) >>> _zz_999);
  assign _zz_8177 = _zz_8178;
  assign _zz_8178 = ($signed(data_mid_113_real) - $signed(_zz_997));
  assign _zz_8179 = _zz_8180;
  assign _zz_8180 = ($signed(_zz_8181) >>> _zz_999);
  assign _zz_8181 = _zz_8182;
  assign _zz_8182 = ($signed(data_mid_113_imag) - $signed(_zz_998));
  assign _zz_8183 = _zz_8184;
  assign _zz_8184 = ($signed(_zz_8185) >>> _zz_1000);
  assign _zz_8185 = _zz_8186;
  assign _zz_8186 = ($signed(data_mid_113_real) + $signed(_zz_997));
  assign _zz_8187 = _zz_8188;
  assign _zz_8188 = ($signed(_zz_8189) >>> _zz_1000);
  assign _zz_8189 = _zz_8190;
  assign _zz_8190 = ($signed(data_mid_113_imag) + $signed(_zz_998));
  assign _zz_8191 = ($signed(twiddle_factor_table_9_real) * $signed(data_mid_122_real));
  assign _zz_8192 = ($signed(twiddle_factor_table_9_imag) * $signed(data_mid_122_imag));
  assign _zz_8193 = fixTo_500_dout;
  assign _zz_8194 = ($signed(twiddle_factor_table_9_real) * $signed(data_mid_122_imag));
  assign _zz_8195 = ($signed(twiddle_factor_table_9_imag) * $signed(data_mid_122_real));
  assign _zz_8196 = fixTo_501_dout;
  assign _zz_8197 = _zz_8198;
  assign _zz_8198 = ($signed(_zz_8199) >>> _zz_1003);
  assign _zz_8199 = _zz_8200;
  assign _zz_8200 = ($signed(data_mid_114_real) - $signed(_zz_1001));
  assign _zz_8201 = _zz_8202;
  assign _zz_8202 = ($signed(_zz_8203) >>> _zz_1003);
  assign _zz_8203 = _zz_8204;
  assign _zz_8204 = ($signed(data_mid_114_imag) - $signed(_zz_1002));
  assign _zz_8205 = _zz_8206;
  assign _zz_8206 = ($signed(_zz_8207) >>> _zz_1004);
  assign _zz_8207 = _zz_8208;
  assign _zz_8208 = ($signed(data_mid_114_real) + $signed(_zz_1001));
  assign _zz_8209 = _zz_8210;
  assign _zz_8210 = ($signed(_zz_8211) >>> _zz_1004);
  assign _zz_8211 = _zz_8212;
  assign _zz_8212 = ($signed(data_mid_114_imag) + $signed(_zz_1002));
  assign _zz_8213 = ($signed(twiddle_factor_table_10_real) * $signed(data_mid_123_real));
  assign _zz_8214 = ($signed(twiddle_factor_table_10_imag) * $signed(data_mid_123_imag));
  assign _zz_8215 = fixTo_502_dout;
  assign _zz_8216 = ($signed(twiddle_factor_table_10_real) * $signed(data_mid_123_imag));
  assign _zz_8217 = ($signed(twiddle_factor_table_10_imag) * $signed(data_mid_123_real));
  assign _zz_8218 = fixTo_503_dout;
  assign _zz_8219 = _zz_8220;
  assign _zz_8220 = ($signed(_zz_8221) >>> _zz_1007);
  assign _zz_8221 = _zz_8222;
  assign _zz_8222 = ($signed(data_mid_115_real) - $signed(_zz_1005));
  assign _zz_8223 = _zz_8224;
  assign _zz_8224 = ($signed(_zz_8225) >>> _zz_1007);
  assign _zz_8225 = _zz_8226;
  assign _zz_8226 = ($signed(data_mid_115_imag) - $signed(_zz_1006));
  assign _zz_8227 = _zz_8228;
  assign _zz_8228 = ($signed(_zz_8229) >>> _zz_1008);
  assign _zz_8229 = _zz_8230;
  assign _zz_8230 = ($signed(data_mid_115_real) + $signed(_zz_1005));
  assign _zz_8231 = _zz_8232;
  assign _zz_8232 = ($signed(_zz_8233) >>> _zz_1008);
  assign _zz_8233 = _zz_8234;
  assign _zz_8234 = ($signed(data_mid_115_imag) + $signed(_zz_1006));
  assign _zz_8235 = ($signed(twiddle_factor_table_11_real) * $signed(data_mid_124_real));
  assign _zz_8236 = ($signed(twiddle_factor_table_11_imag) * $signed(data_mid_124_imag));
  assign _zz_8237 = fixTo_504_dout;
  assign _zz_8238 = ($signed(twiddle_factor_table_11_real) * $signed(data_mid_124_imag));
  assign _zz_8239 = ($signed(twiddle_factor_table_11_imag) * $signed(data_mid_124_real));
  assign _zz_8240 = fixTo_505_dout;
  assign _zz_8241 = _zz_8242;
  assign _zz_8242 = ($signed(_zz_8243) >>> _zz_1011);
  assign _zz_8243 = _zz_8244;
  assign _zz_8244 = ($signed(data_mid_116_real) - $signed(_zz_1009));
  assign _zz_8245 = _zz_8246;
  assign _zz_8246 = ($signed(_zz_8247) >>> _zz_1011);
  assign _zz_8247 = _zz_8248;
  assign _zz_8248 = ($signed(data_mid_116_imag) - $signed(_zz_1010));
  assign _zz_8249 = _zz_8250;
  assign _zz_8250 = ($signed(_zz_8251) >>> _zz_1012);
  assign _zz_8251 = _zz_8252;
  assign _zz_8252 = ($signed(data_mid_116_real) + $signed(_zz_1009));
  assign _zz_8253 = _zz_8254;
  assign _zz_8254 = ($signed(_zz_8255) >>> _zz_1012);
  assign _zz_8255 = _zz_8256;
  assign _zz_8256 = ($signed(data_mid_116_imag) + $signed(_zz_1010));
  assign _zz_8257 = ($signed(twiddle_factor_table_12_real) * $signed(data_mid_125_real));
  assign _zz_8258 = ($signed(twiddle_factor_table_12_imag) * $signed(data_mid_125_imag));
  assign _zz_8259 = fixTo_506_dout;
  assign _zz_8260 = ($signed(twiddle_factor_table_12_real) * $signed(data_mid_125_imag));
  assign _zz_8261 = ($signed(twiddle_factor_table_12_imag) * $signed(data_mid_125_real));
  assign _zz_8262 = fixTo_507_dout;
  assign _zz_8263 = _zz_8264;
  assign _zz_8264 = ($signed(_zz_8265) >>> _zz_1015);
  assign _zz_8265 = _zz_8266;
  assign _zz_8266 = ($signed(data_mid_117_real) - $signed(_zz_1013));
  assign _zz_8267 = _zz_8268;
  assign _zz_8268 = ($signed(_zz_8269) >>> _zz_1015);
  assign _zz_8269 = _zz_8270;
  assign _zz_8270 = ($signed(data_mid_117_imag) - $signed(_zz_1014));
  assign _zz_8271 = _zz_8272;
  assign _zz_8272 = ($signed(_zz_8273) >>> _zz_1016);
  assign _zz_8273 = _zz_8274;
  assign _zz_8274 = ($signed(data_mid_117_real) + $signed(_zz_1013));
  assign _zz_8275 = _zz_8276;
  assign _zz_8276 = ($signed(_zz_8277) >>> _zz_1016);
  assign _zz_8277 = _zz_8278;
  assign _zz_8278 = ($signed(data_mid_117_imag) + $signed(_zz_1014));
  assign _zz_8279 = ($signed(twiddle_factor_table_13_real) * $signed(data_mid_126_real));
  assign _zz_8280 = ($signed(twiddle_factor_table_13_imag) * $signed(data_mid_126_imag));
  assign _zz_8281 = fixTo_508_dout;
  assign _zz_8282 = ($signed(twiddle_factor_table_13_real) * $signed(data_mid_126_imag));
  assign _zz_8283 = ($signed(twiddle_factor_table_13_imag) * $signed(data_mid_126_real));
  assign _zz_8284 = fixTo_509_dout;
  assign _zz_8285 = _zz_8286;
  assign _zz_8286 = ($signed(_zz_8287) >>> _zz_1019);
  assign _zz_8287 = _zz_8288;
  assign _zz_8288 = ($signed(data_mid_118_real) - $signed(_zz_1017));
  assign _zz_8289 = _zz_8290;
  assign _zz_8290 = ($signed(_zz_8291) >>> _zz_1019);
  assign _zz_8291 = _zz_8292;
  assign _zz_8292 = ($signed(data_mid_118_imag) - $signed(_zz_1018));
  assign _zz_8293 = _zz_8294;
  assign _zz_8294 = ($signed(_zz_8295) >>> _zz_1020);
  assign _zz_8295 = _zz_8296;
  assign _zz_8296 = ($signed(data_mid_118_real) + $signed(_zz_1017));
  assign _zz_8297 = _zz_8298;
  assign _zz_8298 = ($signed(_zz_8299) >>> _zz_1020);
  assign _zz_8299 = _zz_8300;
  assign _zz_8300 = ($signed(data_mid_118_imag) + $signed(_zz_1018));
  assign _zz_8301 = ($signed(twiddle_factor_table_14_real) * $signed(data_mid_127_real));
  assign _zz_8302 = ($signed(twiddle_factor_table_14_imag) * $signed(data_mid_127_imag));
  assign _zz_8303 = fixTo_510_dout;
  assign _zz_8304 = ($signed(twiddle_factor_table_14_real) * $signed(data_mid_127_imag));
  assign _zz_8305 = ($signed(twiddle_factor_table_14_imag) * $signed(data_mid_127_real));
  assign _zz_8306 = fixTo_511_dout;
  assign _zz_8307 = _zz_8308;
  assign _zz_8308 = ($signed(_zz_8309) >>> _zz_1023);
  assign _zz_8309 = _zz_8310;
  assign _zz_8310 = ($signed(data_mid_119_real) - $signed(_zz_1021));
  assign _zz_8311 = _zz_8312;
  assign _zz_8312 = ($signed(_zz_8313) >>> _zz_1023);
  assign _zz_8313 = _zz_8314;
  assign _zz_8314 = ($signed(data_mid_119_imag) - $signed(_zz_1022));
  assign _zz_8315 = _zz_8316;
  assign _zz_8316 = ($signed(_zz_8317) >>> _zz_1024);
  assign _zz_8317 = _zz_8318;
  assign _zz_8318 = ($signed(data_mid_119_real) + $signed(_zz_1021));
  assign _zz_8319 = _zz_8320;
  assign _zz_8320 = ($signed(_zz_8321) >>> _zz_1024);
  assign _zz_8321 = _zz_8322;
  assign _zz_8322 = ($signed(data_mid_119_imag) + $signed(_zz_1022));
  assign _zz_8323 = ($signed(twiddle_factor_table_15_real) * $signed(data_mid_16_real));
  assign _zz_8324 = ($signed(twiddle_factor_table_15_imag) * $signed(data_mid_16_imag));
  assign _zz_8325 = fixTo_512_dout;
  assign _zz_8326 = ($signed(twiddle_factor_table_15_real) * $signed(data_mid_16_imag));
  assign _zz_8327 = ($signed(twiddle_factor_table_15_imag) * $signed(data_mid_16_real));
  assign _zz_8328 = fixTo_513_dout;
  assign _zz_8329 = _zz_8330;
  assign _zz_8330 = ($signed(_zz_8331) >>> _zz_1027);
  assign _zz_8331 = _zz_8332;
  assign _zz_8332 = ($signed(data_mid_0_real) - $signed(_zz_1025));
  assign _zz_8333 = _zz_8334;
  assign _zz_8334 = ($signed(_zz_8335) >>> _zz_1027);
  assign _zz_8335 = _zz_8336;
  assign _zz_8336 = ($signed(data_mid_0_imag) - $signed(_zz_1026));
  assign _zz_8337 = _zz_8338;
  assign _zz_8338 = ($signed(_zz_8339) >>> _zz_1028);
  assign _zz_8339 = _zz_8340;
  assign _zz_8340 = ($signed(data_mid_0_real) + $signed(_zz_1025));
  assign _zz_8341 = _zz_8342;
  assign _zz_8342 = ($signed(_zz_8343) >>> _zz_1028);
  assign _zz_8343 = _zz_8344;
  assign _zz_8344 = ($signed(data_mid_0_imag) + $signed(_zz_1026));
  assign _zz_8345 = ($signed(twiddle_factor_table_16_real) * $signed(data_mid_17_real));
  assign _zz_8346 = ($signed(twiddle_factor_table_16_imag) * $signed(data_mid_17_imag));
  assign _zz_8347 = fixTo_514_dout;
  assign _zz_8348 = ($signed(twiddle_factor_table_16_real) * $signed(data_mid_17_imag));
  assign _zz_8349 = ($signed(twiddle_factor_table_16_imag) * $signed(data_mid_17_real));
  assign _zz_8350 = fixTo_515_dout;
  assign _zz_8351 = _zz_8352;
  assign _zz_8352 = ($signed(_zz_8353) >>> _zz_1031);
  assign _zz_8353 = _zz_8354;
  assign _zz_8354 = ($signed(data_mid_1_real) - $signed(_zz_1029));
  assign _zz_8355 = _zz_8356;
  assign _zz_8356 = ($signed(_zz_8357) >>> _zz_1031);
  assign _zz_8357 = _zz_8358;
  assign _zz_8358 = ($signed(data_mid_1_imag) - $signed(_zz_1030));
  assign _zz_8359 = _zz_8360;
  assign _zz_8360 = ($signed(_zz_8361) >>> _zz_1032);
  assign _zz_8361 = _zz_8362;
  assign _zz_8362 = ($signed(data_mid_1_real) + $signed(_zz_1029));
  assign _zz_8363 = _zz_8364;
  assign _zz_8364 = ($signed(_zz_8365) >>> _zz_1032);
  assign _zz_8365 = _zz_8366;
  assign _zz_8366 = ($signed(data_mid_1_imag) + $signed(_zz_1030));
  assign _zz_8367 = ($signed(twiddle_factor_table_17_real) * $signed(data_mid_18_real));
  assign _zz_8368 = ($signed(twiddle_factor_table_17_imag) * $signed(data_mid_18_imag));
  assign _zz_8369 = fixTo_516_dout;
  assign _zz_8370 = ($signed(twiddle_factor_table_17_real) * $signed(data_mid_18_imag));
  assign _zz_8371 = ($signed(twiddle_factor_table_17_imag) * $signed(data_mid_18_real));
  assign _zz_8372 = fixTo_517_dout;
  assign _zz_8373 = _zz_8374;
  assign _zz_8374 = ($signed(_zz_8375) >>> _zz_1035);
  assign _zz_8375 = _zz_8376;
  assign _zz_8376 = ($signed(data_mid_2_real) - $signed(_zz_1033));
  assign _zz_8377 = _zz_8378;
  assign _zz_8378 = ($signed(_zz_8379) >>> _zz_1035);
  assign _zz_8379 = _zz_8380;
  assign _zz_8380 = ($signed(data_mid_2_imag) - $signed(_zz_1034));
  assign _zz_8381 = _zz_8382;
  assign _zz_8382 = ($signed(_zz_8383) >>> _zz_1036);
  assign _zz_8383 = _zz_8384;
  assign _zz_8384 = ($signed(data_mid_2_real) + $signed(_zz_1033));
  assign _zz_8385 = _zz_8386;
  assign _zz_8386 = ($signed(_zz_8387) >>> _zz_1036);
  assign _zz_8387 = _zz_8388;
  assign _zz_8388 = ($signed(data_mid_2_imag) + $signed(_zz_1034));
  assign _zz_8389 = ($signed(twiddle_factor_table_18_real) * $signed(data_mid_19_real));
  assign _zz_8390 = ($signed(twiddle_factor_table_18_imag) * $signed(data_mid_19_imag));
  assign _zz_8391 = fixTo_518_dout;
  assign _zz_8392 = ($signed(twiddle_factor_table_18_real) * $signed(data_mid_19_imag));
  assign _zz_8393 = ($signed(twiddle_factor_table_18_imag) * $signed(data_mid_19_real));
  assign _zz_8394 = fixTo_519_dout;
  assign _zz_8395 = _zz_8396;
  assign _zz_8396 = ($signed(_zz_8397) >>> _zz_1039);
  assign _zz_8397 = _zz_8398;
  assign _zz_8398 = ($signed(data_mid_3_real) - $signed(_zz_1037));
  assign _zz_8399 = _zz_8400;
  assign _zz_8400 = ($signed(_zz_8401) >>> _zz_1039);
  assign _zz_8401 = _zz_8402;
  assign _zz_8402 = ($signed(data_mid_3_imag) - $signed(_zz_1038));
  assign _zz_8403 = _zz_8404;
  assign _zz_8404 = ($signed(_zz_8405) >>> _zz_1040);
  assign _zz_8405 = _zz_8406;
  assign _zz_8406 = ($signed(data_mid_3_real) + $signed(_zz_1037));
  assign _zz_8407 = _zz_8408;
  assign _zz_8408 = ($signed(_zz_8409) >>> _zz_1040);
  assign _zz_8409 = _zz_8410;
  assign _zz_8410 = ($signed(data_mid_3_imag) + $signed(_zz_1038));
  assign _zz_8411 = ($signed(twiddle_factor_table_19_real) * $signed(data_mid_20_real));
  assign _zz_8412 = ($signed(twiddle_factor_table_19_imag) * $signed(data_mid_20_imag));
  assign _zz_8413 = fixTo_520_dout;
  assign _zz_8414 = ($signed(twiddle_factor_table_19_real) * $signed(data_mid_20_imag));
  assign _zz_8415 = ($signed(twiddle_factor_table_19_imag) * $signed(data_mid_20_real));
  assign _zz_8416 = fixTo_521_dout;
  assign _zz_8417 = _zz_8418;
  assign _zz_8418 = ($signed(_zz_8419) >>> _zz_1043);
  assign _zz_8419 = _zz_8420;
  assign _zz_8420 = ($signed(data_mid_4_real) - $signed(_zz_1041));
  assign _zz_8421 = _zz_8422;
  assign _zz_8422 = ($signed(_zz_8423) >>> _zz_1043);
  assign _zz_8423 = _zz_8424;
  assign _zz_8424 = ($signed(data_mid_4_imag) - $signed(_zz_1042));
  assign _zz_8425 = _zz_8426;
  assign _zz_8426 = ($signed(_zz_8427) >>> _zz_1044);
  assign _zz_8427 = _zz_8428;
  assign _zz_8428 = ($signed(data_mid_4_real) + $signed(_zz_1041));
  assign _zz_8429 = _zz_8430;
  assign _zz_8430 = ($signed(_zz_8431) >>> _zz_1044);
  assign _zz_8431 = _zz_8432;
  assign _zz_8432 = ($signed(data_mid_4_imag) + $signed(_zz_1042));
  assign _zz_8433 = ($signed(twiddle_factor_table_20_real) * $signed(data_mid_21_real));
  assign _zz_8434 = ($signed(twiddle_factor_table_20_imag) * $signed(data_mid_21_imag));
  assign _zz_8435 = fixTo_522_dout;
  assign _zz_8436 = ($signed(twiddle_factor_table_20_real) * $signed(data_mid_21_imag));
  assign _zz_8437 = ($signed(twiddle_factor_table_20_imag) * $signed(data_mid_21_real));
  assign _zz_8438 = fixTo_523_dout;
  assign _zz_8439 = _zz_8440;
  assign _zz_8440 = ($signed(_zz_8441) >>> _zz_1047);
  assign _zz_8441 = _zz_8442;
  assign _zz_8442 = ($signed(data_mid_5_real) - $signed(_zz_1045));
  assign _zz_8443 = _zz_8444;
  assign _zz_8444 = ($signed(_zz_8445) >>> _zz_1047);
  assign _zz_8445 = _zz_8446;
  assign _zz_8446 = ($signed(data_mid_5_imag) - $signed(_zz_1046));
  assign _zz_8447 = _zz_8448;
  assign _zz_8448 = ($signed(_zz_8449) >>> _zz_1048);
  assign _zz_8449 = _zz_8450;
  assign _zz_8450 = ($signed(data_mid_5_real) + $signed(_zz_1045));
  assign _zz_8451 = _zz_8452;
  assign _zz_8452 = ($signed(_zz_8453) >>> _zz_1048);
  assign _zz_8453 = _zz_8454;
  assign _zz_8454 = ($signed(data_mid_5_imag) + $signed(_zz_1046));
  assign _zz_8455 = ($signed(twiddle_factor_table_21_real) * $signed(data_mid_22_real));
  assign _zz_8456 = ($signed(twiddle_factor_table_21_imag) * $signed(data_mid_22_imag));
  assign _zz_8457 = fixTo_524_dout;
  assign _zz_8458 = ($signed(twiddle_factor_table_21_real) * $signed(data_mid_22_imag));
  assign _zz_8459 = ($signed(twiddle_factor_table_21_imag) * $signed(data_mid_22_real));
  assign _zz_8460 = fixTo_525_dout;
  assign _zz_8461 = _zz_8462;
  assign _zz_8462 = ($signed(_zz_8463) >>> _zz_1051);
  assign _zz_8463 = _zz_8464;
  assign _zz_8464 = ($signed(data_mid_6_real) - $signed(_zz_1049));
  assign _zz_8465 = _zz_8466;
  assign _zz_8466 = ($signed(_zz_8467) >>> _zz_1051);
  assign _zz_8467 = _zz_8468;
  assign _zz_8468 = ($signed(data_mid_6_imag) - $signed(_zz_1050));
  assign _zz_8469 = _zz_8470;
  assign _zz_8470 = ($signed(_zz_8471) >>> _zz_1052);
  assign _zz_8471 = _zz_8472;
  assign _zz_8472 = ($signed(data_mid_6_real) + $signed(_zz_1049));
  assign _zz_8473 = _zz_8474;
  assign _zz_8474 = ($signed(_zz_8475) >>> _zz_1052);
  assign _zz_8475 = _zz_8476;
  assign _zz_8476 = ($signed(data_mid_6_imag) + $signed(_zz_1050));
  assign _zz_8477 = ($signed(twiddle_factor_table_22_real) * $signed(data_mid_23_real));
  assign _zz_8478 = ($signed(twiddle_factor_table_22_imag) * $signed(data_mid_23_imag));
  assign _zz_8479 = fixTo_526_dout;
  assign _zz_8480 = ($signed(twiddle_factor_table_22_real) * $signed(data_mid_23_imag));
  assign _zz_8481 = ($signed(twiddle_factor_table_22_imag) * $signed(data_mid_23_real));
  assign _zz_8482 = fixTo_527_dout;
  assign _zz_8483 = _zz_8484;
  assign _zz_8484 = ($signed(_zz_8485) >>> _zz_1055);
  assign _zz_8485 = _zz_8486;
  assign _zz_8486 = ($signed(data_mid_7_real) - $signed(_zz_1053));
  assign _zz_8487 = _zz_8488;
  assign _zz_8488 = ($signed(_zz_8489) >>> _zz_1055);
  assign _zz_8489 = _zz_8490;
  assign _zz_8490 = ($signed(data_mid_7_imag) - $signed(_zz_1054));
  assign _zz_8491 = _zz_8492;
  assign _zz_8492 = ($signed(_zz_8493) >>> _zz_1056);
  assign _zz_8493 = _zz_8494;
  assign _zz_8494 = ($signed(data_mid_7_real) + $signed(_zz_1053));
  assign _zz_8495 = _zz_8496;
  assign _zz_8496 = ($signed(_zz_8497) >>> _zz_1056);
  assign _zz_8497 = _zz_8498;
  assign _zz_8498 = ($signed(data_mid_7_imag) + $signed(_zz_1054));
  assign _zz_8499 = ($signed(twiddle_factor_table_23_real) * $signed(data_mid_24_real));
  assign _zz_8500 = ($signed(twiddle_factor_table_23_imag) * $signed(data_mid_24_imag));
  assign _zz_8501 = fixTo_528_dout;
  assign _zz_8502 = ($signed(twiddle_factor_table_23_real) * $signed(data_mid_24_imag));
  assign _zz_8503 = ($signed(twiddle_factor_table_23_imag) * $signed(data_mid_24_real));
  assign _zz_8504 = fixTo_529_dout;
  assign _zz_8505 = _zz_8506;
  assign _zz_8506 = ($signed(_zz_8507) >>> _zz_1059);
  assign _zz_8507 = _zz_8508;
  assign _zz_8508 = ($signed(data_mid_8_real) - $signed(_zz_1057));
  assign _zz_8509 = _zz_8510;
  assign _zz_8510 = ($signed(_zz_8511) >>> _zz_1059);
  assign _zz_8511 = _zz_8512;
  assign _zz_8512 = ($signed(data_mid_8_imag) - $signed(_zz_1058));
  assign _zz_8513 = _zz_8514;
  assign _zz_8514 = ($signed(_zz_8515) >>> _zz_1060);
  assign _zz_8515 = _zz_8516;
  assign _zz_8516 = ($signed(data_mid_8_real) + $signed(_zz_1057));
  assign _zz_8517 = _zz_8518;
  assign _zz_8518 = ($signed(_zz_8519) >>> _zz_1060);
  assign _zz_8519 = _zz_8520;
  assign _zz_8520 = ($signed(data_mid_8_imag) + $signed(_zz_1058));
  assign _zz_8521 = ($signed(twiddle_factor_table_24_real) * $signed(data_mid_25_real));
  assign _zz_8522 = ($signed(twiddle_factor_table_24_imag) * $signed(data_mid_25_imag));
  assign _zz_8523 = fixTo_530_dout;
  assign _zz_8524 = ($signed(twiddle_factor_table_24_real) * $signed(data_mid_25_imag));
  assign _zz_8525 = ($signed(twiddle_factor_table_24_imag) * $signed(data_mid_25_real));
  assign _zz_8526 = fixTo_531_dout;
  assign _zz_8527 = _zz_8528;
  assign _zz_8528 = ($signed(_zz_8529) >>> _zz_1063);
  assign _zz_8529 = _zz_8530;
  assign _zz_8530 = ($signed(data_mid_9_real) - $signed(_zz_1061));
  assign _zz_8531 = _zz_8532;
  assign _zz_8532 = ($signed(_zz_8533) >>> _zz_1063);
  assign _zz_8533 = _zz_8534;
  assign _zz_8534 = ($signed(data_mid_9_imag) - $signed(_zz_1062));
  assign _zz_8535 = _zz_8536;
  assign _zz_8536 = ($signed(_zz_8537) >>> _zz_1064);
  assign _zz_8537 = _zz_8538;
  assign _zz_8538 = ($signed(data_mid_9_real) + $signed(_zz_1061));
  assign _zz_8539 = _zz_8540;
  assign _zz_8540 = ($signed(_zz_8541) >>> _zz_1064);
  assign _zz_8541 = _zz_8542;
  assign _zz_8542 = ($signed(data_mid_9_imag) + $signed(_zz_1062));
  assign _zz_8543 = ($signed(twiddle_factor_table_25_real) * $signed(data_mid_26_real));
  assign _zz_8544 = ($signed(twiddle_factor_table_25_imag) * $signed(data_mid_26_imag));
  assign _zz_8545 = fixTo_532_dout;
  assign _zz_8546 = ($signed(twiddle_factor_table_25_real) * $signed(data_mid_26_imag));
  assign _zz_8547 = ($signed(twiddle_factor_table_25_imag) * $signed(data_mid_26_real));
  assign _zz_8548 = fixTo_533_dout;
  assign _zz_8549 = _zz_8550;
  assign _zz_8550 = ($signed(_zz_8551) >>> _zz_1067);
  assign _zz_8551 = _zz_8552;
  assign _zz_8552 = ($signed(data_mid_10_real) - $signed(_zz_1065));
  assign _zz_8553 = _zz_8554;
  assign _zz_8554 = ($signed(_zz_8555) >>> _zz_1067);
  assign _zz_8555 = _zz_8556;
  assign _zz_8556 = ($signed(data_mid_10_imag) - $signed(_zz_1066));
  assign _zz_8557 = _zz_8558;
  assign _zz_8558 = ($signed(_zz_8559) >>> _zz_1068);
  assign _zz_8559 = _zz_8560;
  assign _zz_8560 = ($signed(data_mid_10_real) + $signed(_zz_1065));
  assign _zz_8561 = _zz_8562;
  assign _zz_8562 = ($signed(_zz_8563) >>> _zz_1068);
  assign _zz_8563 = _zz_8564;
  assign _zz_8564 = ($signed(data_mid_10_imag) + $signed(_zz_1066));
  assign _zz_8565 = ($signed(twiddle_factor_table_26_real) * $signed(data_mid_27_real));
  assign _zz_8566 = ($signed(twiddle_factor_table_26_imag) * $signed(data_mid_27_imag));
  assign _zz_8567 = fixTo_534_dout;
  assign _zz_8568 = ($signed(twiddle_factor_table_26_real) * $signed(data_mid_27_imag));
  assign _zz_8569 = ($signed(twiddle_factor_table_26_imag) * $signed(data_mid_27_real));
  assign _zz_8570 = fixTo_535_dout;
  assign _zz_8571 = _zz_8572;
  assign _zz_8572 = ($signed(_zz_8573) >>> _zz_1071);
  assign _zz_8573 = _zz_8574;
  assign _zz_8574 = ($signed(data_mid_11_real) - $signed(_zz_1069));
  assign _zz_8575 = _zz_8576;
  assign _zz_8576 = ($signed(_zz_8577) >>> _zz_1071);
  assign _zz_8577 = _zz_8578;
  assign _zz_8578 = ($signed(data_mid_11_imag) - $signed(_zz_1070));
  assign _zz_8579 = _zz_8580;
  assign _zz_8580 = ($signed(_zz_8581) >>> _zz_1072);
  assign _zz_8581 = _zz_8582;
  assign _zz_8582 = ($signed(data_mid_11_real) + $signed(_zz_1069));
  assign _zz_8583 = _zz_8584;
  assign _zz_8584 = ($signed(_zz_8585) >>> _zz_1072);
  assign _zz_8585 = _zz_8586;
  assign _zz_8586 = ($signed(data_mid_11_imag) + $signed(_zz_1070));
  assign _zz_8587 = ($signed(twiddle_factor_table_27_real) * $signed(data_mid_28_real));
  assign _zz_8588 = ($signed(twiddle_factor_table_27_imag) * $signed(data_mid_28_imag));
  assign _zz_8589 = fixTo_536_dout;
  assign _zz_8590 = ($signed(twiddle_factor_table_27_real) * $signed(data_mid_28_imag));
  assign _zz_8591 = ($signed(twiddle_factor_table_27_imag) * $signed(data_mid_28_real));
  assign _zz_8592 = fixTo_537_dout;
  assign _zz_8593 = _zz_8594;
  assign _zz_8594 = ($signed(_zz_8595) >>> _zz_1075);
  assign _zz_8595 = _zz_8596;
  assign _zz_8596 = ($signed(data_mid_12_real) - $signed(_zz_1073));
  assign _zz_8597 = _zz_8598;
  assign _zz_8598 = ($signed(_zz_8599) >>> _zz_1075);
  assign _zz_8599 = _zz_8600;
  assign _zz_8600 = ($signed(data_mid_12_imag) - $signed(_zz_1074));
  assign _zz_8601 = _zz_8602;
  assign _zz_8602 = ($signed(_zz_8603) >>> _zz_1076);
  assign _zz_8603 = _zz_8604;
  assign _zz_8604 = ($signed(data_mid_12_real) + $signed(_zz_1073));
  assign _zz_8605 = _zz_8606;
  assign _zz_8606 = ($signed(_zz_8607) >>> _zz_1076);
  assign _zz_8607 = _zz_8608;
  assign _zz_8608 = ($signed(data_mid_12_imag) + $signed(_zz_1074));
  assign _zz_8609 = ($signed(twiddle_factor_table_28_real) * $signed(data_mid_29_real));
  assign _zz_8610 = ($signed(twiddle_factor_table_28_imag) * $signed(data_mid_29_imag));
  assign _zz_8611 = fixTo_538_dout;
  assign _zz_8612 = ($signed(twiddle_factor_table_28_real) * $signed(data_mid_29_imag));
  assign _zz_8613 = ($signed(twiddle_factor_table_28_imag) * $signed(data_mid_29_real));
  assign _zz_8614 = fixTo_539_dout;
  assign _zz_8615 = _zz_8616;
  assign _zz_8616 = ($signed(_zz_8617) >>> _zz_1079);
  assign _zz_8617 = _zz_8618;
  assign _zz_8618 = ($signed(data_mid_13_real) - $signed(_zz_1077));
  assign _zz_8619 = _zz_8620;
  assign _zz_8620 = ($signed(_zz_8621) >>> _zz_1079);
  assign _zz_8621 = _zz_8622;
  assign _zz_8622 = ($signed(data_mid_13_imag) - $signed(_zz_1078));
  assign _zz_8623 = _zz_8624;
  assign _zz_8624 = ($signed(_zz_8625) >>> _zz_1080);
  assign _zz_8625 = _zz_8626;
  assign _zz_8626 = ($signed(data_mid_13_real) + $signed(_zz_1077));
  assign _zz_8627 = _zz_8628;
  assign _zz_8628 = ($signed(_zz_8629) >>> _zz_1080);
  assign _zz_8629 = _zz_8630;
  assign _zz_8630 = ($signed(data_mid_13_imag) + $signed(_zz_1078));
  assign _zz_8631 = ($signed(twiddle_factor_table_29_real) * $signed(data_mid_30_real));
  assign _zz_8632 = ($signed(twiddle_factor_table_29_imag) * $signed(data_mid_30_imag));
  assign _zz_8633 = fixTo_540_dout;
  assign _zz_8634 = ($signed(twiddle_factor_table_29_real) * $signed(data_mid_30_imag));
  assign _zz_8635 = ($signed(twiddle_factor_table_29_imag) * $signed(data_mid_30_real));
  assign _zz_8636 = fixTo_541_dout;
  assign _zz_8637 = _zz_8638;
  assign _zz_8638 = ($signed(_zz_8639) >>> _zz_1083);
  assign _zz_8639 = _zz_8640;
  assign _zz_8640 = ($signed(data_mid_14_real) - $signed(_zz_1081));
  assign _zz_8641 = _zz_8642;
  assign _zz_8642 = ($signed(_zz_8643) >>> _zz_1083);
  assign _zz_8643 = _zz_8644;
  assign _zz_8644 = ($signed(data_mid_14_imag) - $signed(_zz_1082));
  assign _zz_8645 = _zz_8646;
  assign _zz_8646 = ($signed(_zz_8647) >>> _zz_1084);
  assign _zz_8647 = _zz_8648;
  assign _zz_8648 = ($signed(data_mid_14_real) + $signed(_zz_1081));
  assign _zz_8649 = _zz_8650;
  assign _zz_8650 = ($signed(_zz_8651) >>> _zz_1084);
  assign _zz_8651 = _zz_8652;
  assign _zz_8652 = ($signed(data_mid_14_imag) + $signed(_zz_1082));
  assign _zz_8653 = ($signed(twiddle_factor_table_30_real) * $signed(data_mid_31_real));
  assign _zz_8654 = ($signed(twiddle_factor_table_30_imag) * $signed(data_mid_31_imag));
  assign _zz_8655 = fixTo_542_dout;
  assign _zz_8656 = ($signed(twiddle_factor_table_30_real) * $signed(data_mid_31_imag));
  assign _zz_8657 = ($signed(twiddle_factor_table_30_imag) * $signed(data_mid_31_real));
  assign _zz_8658 = fixTo_543_dout;
  assign _zz_8659 = _zz_8660;
  assign _zz_8660 = ($signed(_zz_8661) >>> _zz_1087);
  assign _zz_8661 = _zz_8662;
  assign _zz_8662 = ($signed(data_mid_15_real) - $signed(_zz_1085));
  assign _zz_8663 = _zz_8664;
  assign _zz_8664 = ($signed(_zz_8665) >>> _zz_1087);
  assign _zz_8665 = _zz_8666;
  assign _zz_8666 = ($signed(data_mid_15_imag) - $signed(_zz_1086));
  assign _zz_8667 = _zz_8668;
  assign _zz_8668 = ($signed(_zz_8669) >>> _zz_1088);
  assign _zz_8669 = _zz_8670;
  assign _zz_8670 = ($signed(data_mid_15_real) + $signed(_zz_1085));
  assign _zz_8671 = _zz_8672;
  assign _zz_8672 = ($signed(_zz_8673) >>> _zz_1088);
  assign _zz_8673 = _zz_8674;
  assign _zz_8674 = ($signed(data_mid_15_imag) + $signed(_zz_1086));
  assign _zz_8675 = ($signed(twiddle_factor_table_15_real) * $signed(data_mid_48_real));
  assign _zz_8676 = ($signed(twiddle_factor_table_15_imag) * $signed(data_mid_48_imag));
  assign _zz_8677 = fixTo_544_dout;
  assign _zz_8678 = ($signed(twiddle_factor_table_15_real) * $signed(data_mid_48_imag));
  assign _zz_8679 = ($signed(twiddle_factor_table_15_imag) * $signed(data_mid_48_real));
  assign _zz_8680 = fixTo_545_dout;
  assign _zz_8681 = _zz_8682;
  assign _zz_8682 = ($signed(_zz_8683) >>> _zz_1091);
  assign _zz_8683 = _zz_8684;
  assign _zz_8684 = ($signed(data_mid_32_real) - $signed(_zz_1089));
  assign _zz_8685 = _zz_8686;
  assign _zz_8686 = ($signed(_zz_8687) >>> _zz_1091);
  assign _zz_8687 = _zz_8688;
  assign _zz_8688 = ($signed(data_mid_32_imag) - $signed(_zz_1090));
  assign _zz_8689 = _zz_8690;
  assign _zz_8690 = ($signed(_zz_8691) >>> _zz_1092);
  assign _zz_8691 = _zz_8692;
  assign _zz_8692 = ($signed(data_mid_32_real) + $signed(_zz_1089));
  assign _zz_8693 = _zz_8694;
  assign _zz_8694 = ($signed(_zz_8695) >>> _zz_1092);
  assign _zz_8695 = _zz_8696;
  assign _zz_8696 = ($signed(data_mid_32_imag) + $signed(_zz_1090));
  assign _zz_8697 = ($signed(twiddle_factor_table_16_real) * $signed(data_mid_49_real));
  assign _zz_8698 = ($signed(twiddle_factor_table_16_imag) * $signed(data_mid_49_imag));
  assign _zz_8699 = fixTo_546_dout;
  assign _zz_8700 = ($signed(twiddle_factor_table_16_real) * $signed(data_mid_49_imag));
  assign _zz_8701 = ($signed(twiddle_factor_table_16_imag) * $signed(data_mid_49_real));
  assign _zz_8702 = fixTo_547_dout;
  assign _zz_8703 = _zz_8704;
  assign _zz_8704 = ($signed(_zz_8705) >>> _zz_1095);
  assign _zz_8705 = _zz_8706;
  assign _zz_8706 = ($signed(data_mid_33_real) - $signed(_zz_1093));
  assign _zz_8707 = _zz_8708;
  assign _zz_8708 = ($signed(_zz_8709) >>> _zz_1095);
  assign _zz_8709 = _zz_8710;
  assign _zz_8710 = ($signed(data_mid_33_imag) - $signed(_zz_1094));
  assign _zz_8711 = _zz_8712;
  assign _zz_8712 = ($signed(_zz_8713) >>> _zz_1096);
  assign _zz_8713 = _zz_8714;
  assign _zz_8714 = ($signed(data_mid_33_real) + $signed(_zz_1093));
  assign _zz_8715 = _zz_8716;
  assign _zz_8716 = ($signed(_zz_8717) >>> _zz_1096);
  assign _zz_8717 = _zz_8718;
  assign _zz_8718 = ($signed(data_mid_33_imag) + $signed(_zz_1094));
  assign _zz_8719 = ($signed(twiddle_factor_table_17_real) * $signed(data_mid_50_real));
  assign _zz_8720 = ($signed(twiddle_factor_table_17_imag) * $signed(data_mid_50_imag));
  assign _zz_8721 = fixTo_548_dout;
  assign _zz_8722 = ($signed(twiddle_factor_table_17_real) * $signed(data_mid_50_imag));
  assign _zz_8723 = ($signed(twiddle_factor_table_17_imag) * $signed(data_mid_50_real));
  assign _zz_8724 = fixTo_549_dout;
  assign _zz_8725 = _zz_8726;
  assign _zz_8726 = ($signed(_zz_8727) >>> _zz_1099);
  assign _zz_8727 = _zz_8728;
  assign _zz_8728 = ($signed(data_mid_34_real) - $signed(_zz_1097));
  assign _zz_8729 = _zz_8730;
  assign _zz_8730 = ($signed(_zz_8731) >>> _zz_1099);
  assign _zz_8731 = _zz_8732;
  assign _zz_8732 = ($signed(data_mid_34_imag) - $signed(_zz_1098));
  assign _zz_8733 = _zz_8734;
  assign _zz_8734 = ($signed(_zz_8735) >>> _zz_1100);
  assign _zz_8735 = _zz_8736;
  assign _zz_8736 = ($signed(data_mid_34_real) + $signed(_zz_1097));
  assign _zz_8737 = _zz_8738;
  assign _zz_8738 = ($signed(_zz_8739) >>> _zz_1100);
  assign _zz_8739 = _zz_8740;
  assign _zz_8740 = ($signed(data_mid_34_imag) + $signed(_zz_1098));
  assign _zz_8741 = ($signed(twiddle_factor_table_18_real) * $signed(data_mid_51_real));
  assign _zz_8742 = ($signed(twiddle_factor_table_18_imag) * $signed(data_mid_51_imag));
  assign _zz_8743 = fixTo_550_dout;
  assign _zz_8744 = ($signed(twiddle_factor_table_18_real) * $signed(data_mid_51_imag));
  assign _zz_8745 = ($signed(twiddle_factor_table_18_imag) * $signed(data_mid_51_real));
  assign _zz_8746 = fixTo_551_dout;
  assign _zz_8747 = _zz_8748;
  assign _zz_8748 = ($signed(_zz_8749) >>> _zz_1103);
  assign _zz_8749 = _zz_8750;
  assign _zz_8750 = ($signed(data_mid_35_real) - $signed(_zz_1101));
  assign _zz_8751 = _zz_8752;
  assign _zz_8752 = ($signed(_zz_8753) >>> _zz_1103);
  assign _zz_8753 = _zz_8754;
  assign _zz_8754 = ($signed(data_mid_35_imag) - $signed(_zz_1102));
  assign _zz_8755 = _zz_8756;
  assign _zz_8756 = ($signed(_zz_8757) >>> _zz_1104);
  assign _zz_8757 = _zz_8758;
  assign _zz_8758 = ($signed(data_mid_35_real) + $signed(_zz_1101));
  assign _zz_8759 = _zz_8760;
  assign _zz_8760 = ($signed(_zz_8761) >>> _zz_1104);
  assign _zz_8761 = _zz_8762;
  assign _zz_8762 = ($signed(data_mid_35_imag) + $signed(_zz_1102));
  assign _zz_8763 = ($signed(twiddle_factor_table_19_real) * $signed(data_mid_52_real));
  assign _zz_8764 = ($signed(twiddle_factor_table_19_imag) * $signed(data_mid_52_imag));
  assign _zz_8765 = fixTo_552_dout;
  assign _zz_8766 = ($signed(twiddle_factor_table_19_real) * $signed(data_mid_52_imag));
  assign _zz_8767 = ($signed(twiddle_factor_table_19_imag) * $signed(data_mid_52_real));
  assign _zz_8768 = fixTo_553_dout;
  assign _zz_8769 = _zz_8770;
  assign _zz_8770 = ($signed(_zz_8771) >>> _zz_1107);
  assign _zz_8771 = _zz_8772;
  assign _zz_8772 = ($signed(data_mid_36_real) - $signed(_zz_1105));
  assign _zz_8773 = _zz_8774;
  assign _zz_8774 = ($signed(_zz_8775) >>> _zz_1107);
  assign _zz_8775 = _zz_8776;
  assign _zz_8776 = ($signed(data_mid_36_imag) - $signed(_zz_1106));
  assign _zz_8777 = _zz_8778;
  assign _zz_8778 = ($signed(_zz_8779) >>> _zz_1108);
  assign _zz_8779 = _zz_8780;
  assign _zz_8780 = ($signed(data_mid_36_real) + $signed(_zz_1105));
  assign _zz_8781 = _zz_8782;
  assign _zz_8782 = ($signed(_zz_8783) >>> _zz_1108);
  assign _zz_8783 = _zz_8784;
  assign _zz_8784 = ($signed(data_mid_36_imag) + $signed(_zz_1106));
  assign _zz_8785 = ($signed(twiddle_factor_table_20_real) * $signed(data_mid_53_real));
  assign _zz_8786 = ($signed(twiddle_factor_table_20_imag) * $signed(data_mid_53_imag));
  assign _zz_8787 = fixTo_554_dout;
  assign _zz_8788 = ($signed(twiddle_factor_table_20_real) * $signed(data_mid_53_imag));
  assign _zz_8789 = ($signed(twiddle_factor_table_20_imag) * $signed(data_mid_53_real));
  assign _zz_8790 = fixTo_555_dout;
  assign _zz_8791 = _zz_8792;
  assign _zz_8792 = ($signed(_zz_8793) >>> _zz_1111);
  assign _zz_8793 = _zz_8794;
  assign _zz_8794 = ($signed(data_mid_37_real) - $signed(_zz_1109));
  assign _zz_8795 = _zz_8796;
  assign _zz_8796 = ($signed(_zz_8797) >>> _zz_1111);
  assign _zz_8797 = _zz_8798;
  assign _zz_8798 = ($signed(data_mid_37_imag) - $signed(_zz_1110));
  assign _zz_8799 = _zz_8800;
  assign _zz_8800 = ($signed(_zz_8801) >>> _zz_1112);
  assign _zz_8801 = _zz_8802;
  assign _zz_8802 = ($signed(data_mid_37_real) + $signed(_zz_1109));
  assign _zz_8803 = _zz_8804;
  assign _zz_8804 = ($signed(_zz_8805) >>> _zz_1112);
  assign _zz_8805 = _zz_8806;
  assign _zz_8806 = ($signed(data_mid_37_imag) + $signed(_zz_1110));
  assign _zz_8807 = ($signed(twiddle_factor_table_21_real) * $signed(data_mid_54_real));
  assign _zz_8808 = ($signed(twiddle_factor_table_21_imag) * $signed(data_mid_54_imag));
  assign _zz_8809 = fixTo_556_dout;
  assign _zz_8810 = ($signed(twiddle_factor_table_21_real) * $signed(data_mid_54_imag));
  assign _zz_8811 = ($signed(twiddle_factor_table_21_imag) * $signed(data_mid_54_real));
  assign _zz_8812 = fixTo_557_dout;
  assign _zz_8813 = _zz_8814;
  assign _zz_8814 = ($signed(_zz_8815) >>> _zz_1115);
  assign _zz_8815 = _zz_8816;
  assign _zz_8816 = ($signed(data_mid_38_real) - $signed(_zz_1113));
  assign _zz_8817 = _zz_8818;
  assign _zz_8818 = ($signed(_zz_8819) >>> _zz_1115);
  assign _zz_8819 = _zz_8820;
  assign _zz_8820 = ($signed(data_mid_38_imag) - $signed(_zz_1114));
  assign _zz_8821 = _zz_8822;
  assign _zz_8822 = ($signed(_zz_8823) >>> _zz_1116);
  assign _zz_8823 = _zz_8824;
  assign _zz_8824 = ($signed(data_mid_38_real) + $signed(_zz_1113));
  assign _zz_8825 = _zz_8826;
  assign _zz_8826 = ($signed(_zz_8827) >>> _zz_1116);
  assign _zz_8827 = _zz_8828;
  assign _zz_8828 = ($signed(data_mid_38_imag) + $signed(_zz_1114));
  assign _zz_8829 = ($signed(twiddle_factor_table_22_real) * $signed(data_mid_55_real));
  assign _zz_8830 = ($signed(twiddle_factor_table_22_imag) * $signed(data_mid_55_imag));
  assign _zz_8831 = fixTo_558_dout;
  assign _zz_8832 = ($signed(twiddle_factor_table_22_real) * $signed(data_mid_55_imag));
  assign _zz_8833 = ($signed(twiddle_factor_table_22_imag) * $signed(data_mid_55_real));
  assign _zz_8834 = fixTo_559_dout;
  assign _zz_8835 = _zz_8836;
  assign _zz_8836 = ($signed(_zz_8837) >>> _zz_1119);
  assign _zz_8837 = _zz_8838;
  assign _zz_8838 = ($signed(data_mid_39_real) - $signed(_zz_1117));
  assign _zz_8839 = _zz_8840;
  assign _zz_8840 = ($signed(_zz_8841) >>> _zz_1119);
  assign _zz_8841 = _zz_8842;
  assign _zz_8842 = ($signed(data_mid_39_imag) - $signed(_zz_1118));
  assign _zz_8843 = _zz_8844;
  assign _zz_8844 = ($signed(_zz_8845) >>> _zz_1120);
  assign _zz_8845 = _zz_8846;
  assign _zz_8846 = ($signed(data_mid_39_real) + $signed(_zz_1117));
  assign _zz_8847 = _zz_8848;
  assign _zz_8848 = ($signed(_zz_8849) >>> _zz_1120);
  assign _zz_8849 = _zz_8850;
  assign _zz_8850 = ($signed(data_mid_39_imag) + $signed(_zz_1118));
  assign _zz_8851 = ($signed(twiddle_factor_table_23_real) * $signed(data_mid_56_real));
  assign _zz_8852 = ($signed(twiddle_factor_table_23_imag) * $signed(data_mid_56_imag));
  assign _zz_8853 = fixTo_560_dout;
  assign _zz_8854 = ($signed(twiddle_factor_table_23_real) * $signed(data_mid_56_imag));
  assign _zz_8855 = ($signed(twiddle_factor_table_23_imag) * $signed(data_mid_56_real));
  assign _zz_8856 = fixTo_561_dout;
  assign _zz_8857 = _zz_8858;
  assign _zz_8858 = ($signed(_zz_8859) >>> _zz_1123);
  assign _zz_8859 = _zz_8860;
  assign _zz_8860 = ($signed(data_mid_40_real) - $signed(_zz_1121));
  assign _zz_8861 = _zz_8862;
  assign _zz_8862 = ($signed(_zz_8863) >>> _zz_1123);
  assign _zz_8863 = _zz_8864;
  assign _zz_8864 = ($signed(data_mid_40_imag) - $signed(_zz_1122));
  assign _zz_8865 = _zz_8866;
  assign _zz_8866 = ($signed(_zz_8867) >>> _zz_1124);
  assign _zz_8867 = _zz_8868;
  assign _zz_8868 = ($signed(data_mid_40_real) + $signed(_zz_1121));
  assign _zz_8869 = _zz_8870;
  assign _zz_8870 = ($signed(_zz_8871) >>> _zz_1124);
  assign _zz_8871 = _zz_8872;
  assign _zz_8872 = ($signed(data_mid_40_imag) + $signed(_zz_1122));
  assign _zz_8873 = ($signed(twiddle_factor_table_24_real) * $signed(data_mid_57_real));
  assign _zz_8874 = ($signed(twiddle_factor_table_24_imag) * $signed(data_mid_57_imag));
  assign _zz_8875 = fixTo_562_dout;
  assign _zz_8876 = ($signed(twiddle_factor_table_24_real) * $signed(data_mid_57_imag));
  assign _zz_8877 = ($signed(twiddle_factor_table_24_imag) * $signed(data_mid_57_real));
  assign _zz_8878 = fixTo_563_dout;
  assign _zz_8879 = _zz_8880;
  assign _zz_8880 = ($signed(_zz_8881) >>> _zz_1127);
  assign _zz_8881 = _zz_8882;
  assign _zz_8882 = ($signed(data_mid_41_real) - $signed(_zz_1125));
  assign _zz_8883 = _zz_8884;
  assign _zz_8884 = ($signed(_zz_8885) >>> _zz_1127);
  assign _zz_8885 = _zz_8886;
  assign _zz_8886 = ($signed(data_mid_41_imag) - $signed(_zz_1126));
  assign _zz_8887 = _zz_8888;
  assign _zz_8888 = ($signed(_zz_8889) >>> _zz_1128);
  assign _zz_8889 = _zz_8890;
  assign _zz_8890 = ($signed(data_mid_41_real) + $signed(_zz_1125));
  assign _zz_8891 = _zz_8892;
  assign _zz_8892 = ($signed(_zz_8893) >>> _zz_1128);
  assign _zz_8893 = _zz_8894;
  assign _zz_8894 = ($signed(data_mid_41_imag) + $signed(_zz_1126));
  assign _zz_8895 = ($signed(twiddle_factor_table_25_real) * $signed(data_mid_58_real));
  assign _zz_8896 = ($signed(twiddle_factor_table_25_imag) * $signed(data_mid_58_imag));
  assign _zz_8897 = fixTo_564_dout;
  assign _zz_8898 = ($signed(twiddle_factor_table_25_real) * $signed(data_mid_58_imag));
  assign _zz_8899 = ($signed(twiddle_factor_table_25_imag) * $signed(data_mid_58_real));
  assign _zz_8900 = fixTo_565_dout;
  assign _zz_8901 = _zz_8902;
  assign _zz_8902 = ($signed(_zz_8903) >>> _zz_1131);
  assign _zz_8903 = _zz_8904;
  assign _zz_8904 = ($signed(data_mid_42_real) - $signed(_zz_1129));
  assign _zz_8905 = _zz_8906;
  assign _zz_8906 = ($signed(_zz_8907) >>> _zz_1131);
  assign _zz_8907 = _zz_8908;
  assign _zz_8908 = ($signed(data_mid_42_imag) - $signed(_zz_1130));
  assign _zz_8909 = _zz_8910;
  assign _zz_8910 = ($signed(_zz_8911) >>> _zz_1132);
  assign _zz_8911 = _zz_8912;
  assign _zz_8912 = ($signed(data_mid_42_real) + $signed(_zz_1129));
  assign _zz_8913 = _zz_8914;
  assign _zz_8914 = ($signed(_zz_8915) >>> _zz_1132);
  assign _zz_8915 = _zz_8916;
  assign _zz_8916 = ($signed(data_mid_42_imag) + $signed(_zz_1130));
  assign _zz_8917 = ($signed(twiddle_factor_table_26_real) * $signed(data_mid_59_real));
  assign _zz_8918 = ($signed(twiddle_factor_table_26_imag) * $signed(data_mid_59_imag));
  assign _zz_8919 = fixTo_566_dout;
  assign _zz_8920 = ($signed(twiddle_factor_table_26_real) * $signed(data_mid_59_imag));
  assign _zz_8921 = ($signed(twiddle_factor_table_26_imag) * $signed(data_mid_59_real));
  assign _zz_8922 = fixTo_567_dout;
  assign _zz_8923 = _zz_8924;
  assign _zz_8924 = ($signed(_zz_8925) >>> _zz_1135);
  assign _zz_8925 = _zz_8926;
  assign _zz_8926 = ($signed(data_mid_43_real) - $signed(_zz_1133));
  assign _zz_8927 = _zz_8928;
  assign _zz_8928 = ($signed(_zz_8929) >>> _zz_1135);
  assign _zz_8929 = _zz_8930;
  assign _zz_8930 = ($signed(data_mid_43_imag) - $signed(_zz_1134));
  assign _zz_8931 = _zz_8932;
  assign _zz_8932 = ($signed(_zz_8933) >>> _zz_1136);
  assign _zz_8933 = _zz_8934;
  assign _zz_8934 = ($signed(data_mid_43_real) + $signed(_zz_1133));
  assign _zz_8935 = _zz_8936;
  assign _zz_8936 = ($signed(_zz_8937) >>> _zz_1136);
  assign _zz_8937 = _zz_8938;
  assign _zz_8938 = ($signed(data_mid_43_imag) + $signed(_zz_1134));
  assign _zz_8939 = ($signed(twiddle_factor_table_27_real) * $signed(data_mid_60_real));
  assign _zz_8940 = ($signed(twiddle_factor_table_27_imag) * $signed(data_mid_60_imag));
  assign _zz_8941 = fixTo_568_dout;
  assign _zz_8942 = ($signed(twiddle_factor_table_27_real) * $signed(data_mid_60_imag));
  assign _zz_8943 = ($signed(twiddle_factor_table_27_imag) * $signed(data_mid_60_real));
  assign _zz_8944 = fixTo_569_dout;
  assign _zz_8945 = _zz_8946;
  assign _zz_8946 = ($signed(_zz_8947) >>> _zz_1139);
  assign _zz_8947 = _zz_8948;
  assign _zz_8948 = ($signed(data_mid_44_real) - $signed(_zz_1137));
  assign _zz_8949 = _zz_8950;
  assign _zz_8950 = ($signed(_zz_8951) >>> _zz_1139);
  assign _zz_8951 = _zz_8952;
  assign _zz_8952 = ($signed(data_mid_44_imag) - $signed(_zz_1138));
  assign _zz_8953 = _zz_8954;
  assign _zz_8954 = ($signed(_zz_8955) >>> _zz_1140);
  assign _zz_8955 = _zz_8956;
  assign _zz_8956 = ($signed(data_mid_44_real) + $signed(_zz_1137));
  assign _zz_8957 = _zz_8958;
  assign _zz_8958 = ($signed(_zz_8959) >>> _zz_1140);
  assign _zz_8959 = _zz_8960;
  assign _zz_8960 = ($signed(data_mid_44_imag) + $signed(_zz_1138));
  assign _zz_8961 = ($signed(twiddle_factor_table_28_real) * $signed(data_mid_61_real));
  assign _zz_8962 = ($signed(twiddle_factor_table_28_imag) * $signed(data_mid_61_imag));
  assign _zz_8963 = fixTo_570_dout;
  assign _zz_8964 = ($signed(twiddle_factor_table_28_real) * $signed(data_mid_61_imag));
  assign _zz_8965 = ($signed(twiddle_factor_table_28_imag) * $signed(data_mid_61_real));
  assign _zz_8966 = fixTo_571_dout;
  assign _zz_8967 = _zz_8968;
  assign _zz_8968 = ($signed(_zz_8969) >>> _zz_1143);
  assign _zz_8969 = _zz_8970;
  assign _zz_8970 = ($signed(data_mid_45_real) - $signed(_zz_1141));
  assign _zz_8971 = _zz_8972;
  assign _zz_8972 = ($signed(_zz_8973) >>> _zz_1143);
  assign _zz_8973 = _zz_8974;
  assign _zz_8974 = ($signed(data_mid_45_imag) - $signed(_zz_1142));
  assign _zz_8975 = _zz_8976;
  assign _zz_8976 = ($signed(_zz_8977) >>> _zz_1144);
  assign _zz_8977 = _zz_8978;
  assign _zz_8978 = ($signed(data_mid_45_real) + $signed(_zz_1141));
  assign _zz_8979 = _zz_8980;
  assign _zz_8980 = ($signed(_zz_8981) >>> _zz_1144);
  assign _zz_8981 = _zz_8982;
  assign _zz_8982 = ($signed(data_mid_45_imag) + $signed(_zz_1142));
  assign _zz_8983 = ($signed(twiddle_factor_table_29_real) * $signed(data_mid_62_real));
  assign _zz_8984 = ($signed(twiddle_factor_table_29_imag) * $signed(data_mid_62_imag));
  assign _zz_8985 = fixTo_572_dout;
  assign _zz_8986 = ($signed(twiddle_factor_table_29_real) * $signed(data_mid_62_imag));
  assign _zz_8987 = ($signed(twiddle_factor_table_29_imag) * $signed(data_mid_62_real));
  assign _zz_8988 = fixTo_573_dout;
  assign _zz_8989 = _zz_8990;
  assign _zz_8990 = ($signed(_zz_8991) >>> _zz_1147);
  assign _zz_8991 = _zz_8992;
  assign _zz_8992 = ($signed(data_mid_46_real) - $signed(_zz_1145));
  assign _zz_8993 = _zz_8994;
  assign _zz_8994 = ($signed(_zz_8995) >>> _zz_1147);
  assign _zz_8995 = _zz_8996;
  assign _zz_8996 = ($signed(data_mid_46_imag) - $signed(_zz_1146));
  assign _zz_8997 = _zz_8998;
  assign _zz_8998 = ($signed(_zz_8999) >>> _zz_1148);
  assign _zz_8999 = _zz_9000;
  assign _zz_9000 = ($signed(data_mid_46_real) + $signed(_zz_1145));
  assign _zz_9001 = _zz_9002;
  assign _zz_9002 = ($signed(_zz_9003) >>> _zz_1148);
  assign _zz_9003 = _zz_9004;
  assign _zz_9004 = ($signed(data_mid_46_imag) + $signed(_zz_1146));
  assign _zz_9005 = ($signed(twiddle_factor_table_30_real) * $signed(data_mid_63_real));
  assign _zz_9006 = ($signed(twiddle_factor_table_30_imag) * $signed(data_mid_63_imag));
  assign _zz_9007 = fixTo_574_dout;
  assign _zz_9008 = ($signed(twiddle_factor_table_30_real) * $signed(data_mid_63_imag));
  assign _zz_9009 = ($signed(twiddle_factor_table_30_imag) * $signed(data_mid_63_real));
  assign _zz_9010 = fixTo_575_dout;
  assign _zz_9011 = _zz_9012;
  assign _zz_9012 = ($signed(_zz_9013) >>> _zz_1151);
  assign _zz_9013 = _zz_9014;
  assign _zz_9014 = ($signed(data_mid_47_real) - $signed(_zz_1149));
  assign _zz_9015 = _zz_9016;
  assign _zz_9016 = ($signed(_zz_9017) >>> _zz_1151);
  assign _zz_9017 = _zz_9018;
  assign _zz_9018 = ($signed(data_mid_47_imag) - $signed(_zz_1150));
  assign _zz_9019 = _zz_9020;
  assign _zz_9020 = ($signed(_zz_9021) >>> _zz_1152);
  assign _zz_9021 = _zz_9022;
  assign _zz_9022 = ($signed(data_mid_47_real) + $signed(_zz_1149));
  assign _zz_9023 = _zz_9024;
  assign _zz_9024 = ($signed(_zz_9025) >>> _zz_1152);
  assign _zz_9025 = _zz_9026;
  assign _zz_9026 = ($signed(data_mid_47_imag) + $signed(_zz_1150));
  assign _zz_9027 = ($signed(twiddle_factor_table_15_real) * $signed(data_mid_80_real));
  assign _zz_9028 = ($signed(twiddle_factor_table_15_imag) * $signed(data_mid_80_imag));
  assign _zz_9029 = fixTo_576_dout;
  assign _zz_9030 = ($signed(twiddle_factor_table_15_real) * $signed(data_mid_80_imag));
  assign _zz_9031 = ($signed(twiddle_factor_table_15_imag) * $signed(data_mid_80_real));
  assign _zz_9032 = fixTo_577_dout;
  assign _zz_9033 = _zz_9034;
  assign _zz_9034 = ($signed(_zz_9035) >>> _zz_1155);
  assign _zz_9035 = _zz_9036;
  assign _zz_9036 = ($signed(data_mid_64_real) - $signed(_zz_1153));
  assign _zz_9037 = _zz_9038;
  assign _zz_9038 = ($signed(_zz_9039) >>> _zz_1155);
  assign _zz_9039 = _zz_9040;
  assign _zz_9040 = ($signed(data_mid_64_imag) - $signed(_zz_1154));
  assign _zz_9041 = _zz_9042;
  assign _zz_9042 = ($signed(_zz_9043) >>> _zz_1156);
  assign _zz_9043 = _zz_9044;
  assign _zz_9044 = ($signed(data_mid_64_real) + $signed(_zz_1153));
  assign _zz_9045 = _zz_9046;
  assign _zz_9046 = ($signed(_zz_9047) >>> _zz_1156);
  assign _zz_9047 = _zz_9048;
  assign _zz_9048 = ($signed(data_mid_64_imag) + $signed(_zz_1154));
  assign _zz_9049 = ($signed(twiddle_factor_table_16_real) * $signed(data_mid_81_real));
  assign _zz_9050 = ($signed(twiddle_factor_table_16_imag) * $signed(data_mid_81_imag));
  assign _zz_9051 = fixTo_578_dout;
  assign _zz_9052 = ($signed(twiddle_factor_table_16_real) * $signed(data_mid_81_imag));
  assign _zz_9053 = ($signed(twiddle_factor_table_16_imag) * $signed(data_mid_81_real));
  assign _zz_9054 = fixTo_579_dout;
  assign _zz_9055 = _zz_9056;
  assign _zz_9056 = ($signed(_zz_9057) >>> _zz_1159);
  assign _zz_9057 = _zz_9058;
  assign _zz_9058 = ($signed(data_mid_65_real) - $signed(_zz_1157));
  assign _zz_9059 = _zz_9060;
  assign _zz_9060 = ($signed(_zz_9061) >>> _zz_1159);
  assign _zz_9061 = _zz_9062;
  assign _zz_9062 = ($signed(data_mid_65_imag) - $signed(_zz_1158));
  assign _zz_9063 = _zz_9064;
  assign _zz_9064 = ($signed(_zz_9065) >>> _zz_1160);
  assign _zz_9065 = _zz_9066;
  assign _zz_9066 = ($signed(data_mid_65_real) + $signed(_zz_1157));
  assign _zz_9067 = _zz_9068;
  assign _zz_9068 = ($signed(_zz_9069) >>> _zz_1160);
  assign _zz_9069 = _zz_9070;
  assign _zz_9070 = ($signed(data_mid_65_imag) + $signed(_zz_1158));
  assign _zz_9071 = ($signed(twiddle_factor_table_17_real) * $signed(data_mid_82_real));
  assign _zz_9072 = ($signed(twiddle_factor_table_17_imag) * $signed(data_mid_82_imag));
  assign _zz_9073 = fixTo_580_dout;
  assign _zz_9074 = ($signed(twiddle_factor_table_17_real) * $signed(data_mid_82_imag));
  assign _zz_9075 = ($signed(twiddle_factor_table_17_imag) * $signed(data_mid_82_real));
  assign _zz_9076 = fixTo_581_dout;
  assign _zz_9077 = _zz_9078;
  assign _zz_9078 = ($signed(_zz_9079) >>> _zz_1163);
  assign _zz_9079 = _zz_9080;
  assign _zz_9080 = ($signed(data_mid_66_real) - $signed(_zz_1161));
  assign _zz_9081 = _zz_9082;
  assign _zz_9082 = ($signed(_zz_9083) >>> _zz_1163);
  assign _zz_9083 = _zz_9084;
  assign _zz_9084 = ($signed(data_mid_66_imag) - $signed(_zz_1162));
  assign _zz_9085 = _zz_9086;
  assign _zz_9086 = ($signed(_zz_9087) >>> _zz_1164);
  assign _zz_9087 = _zz_9088;
  assign _zz_9088 = ($signed(data_mid_66_real) + $signed(_zz_1161));
  assign _zz_9089 = _zz_9090;
  assign _zz_9090 = ($signed(_zz_9091) >>> _zz_1164);
  assign _zz_9091 = _zz_9092;
  assign _zz_9092 = ($signed(data_mid_66_imag) + $signed(_zz_1162));
  assign _zz_9093 = ($signed(twiddle_factor_table_18_real) * $signed(data_mid_83_real));
  assign _zz_9094 = ($signed(twiddle_factor_table_18_imag) * $signed(data_mid_83_imag));
  assign _zz_9095 = fixTo_582_dout;
  assign _zz_9096 = ($signed(twiddle_factor_table_18_real) * $signed(data_mid_83_imag));
  assign _zz_9097 = ($signed(twiddle_factor_table_18_imag) * $signed(data_mid_83_real));
  assign _zz_9098 = fixTo_583_dout;
  assign _zz_9099 = _zz_9100;
  assign _zz_9100 = ($signed(_zz_9101) >>> _zz_1167);
  assign _zz_9101 = _zz_9102;
  assign _zz_9102 = ($signed(data_mid_67_real) - $signed(_zz_1165));
  assign _zz_9103 = _zz_9104;
  assign _zz_9104 = ($signed(_zz_9105) >>> _zz_1167);
  assign _zz_9105 = _zz_9106;
  assign _zz_9106 = ($signed(data_mid_67_imag) - $signed(_zz_1166));
  assign _zz_9107 = _zz_9108;
  assign _zz_9108 = ($signed(_zz_9109) >>> _zz_1168);
  assign _zz_9109 = _zz_9110;
  assign _zz_9110 = ($signed(data_mid_67_real) + $signed(_zz_1165));
  assign _zz_9111 = _zz_9112;
  assign _zz_9112 = ($signed(_zz_9113) >>> _zz_1168);
  assign _zz_9113 = _zz_9114;
  assign _zz_9114 = ($signed(data_mid_67_imag) + $signed(_zz_1166));
  assign _zz_9115 = ($signed(twiddle_factor_table_19_real) * $signed(data_mid_84_real));
  assign _zz_9116 = ($signed(twiddle_factor_table_19_imag) * $signed(data_mid_84_imag));
  assign _zz_9117 = fixTo_584_dout;
  assign _zz_9118 = ($signed(twiddle_factor_table_19_real) * $signed(data_mid_84_imag));
  assign _zz_9119 = ($signed(twiddle_factor_table_19_imag) * $signed(data_mid_84_real));
  assign _zz_9120 = fixTo_585_dout;
  assign _zz_9121 = _zz_9122;
  assign _zz_9122 = ($signed(_zz_9123) >>> _zz_1171);
  assign _zz_9123 = _zz_9124;
  assign _zz_9124 = ($signed(data_mid_68_real) - $signed(_zz_1169));
  assign _zz_9125 = _zz_9126;
  assign _zz_9126 = ($signed(_zz_9127) >>> _zz_1171);
  assign _zz_9127 = _zz_9128;
  assign _zz_9128 = ($signed(data_mid_68_imag) - $signed(_zz_1170));
  assign _zz_9129 = _zz_9130;
  assign _zz_9130 = ($signed(_zz_9131) >>> _zz_1172);
  assign _zz_9131 = _zz_9132;
  assign _zz_9132 = ($signed(data_mid_68_real) + $signed(_zz_1169));
  assign _zz_9133 = _zz_9134;
  assign _zz_9134 = ($signed(_zz_9135) >>> _zz_1172);
  assign _zz_9135 = _zz_9136;
  assign _zz_9136 = ($signed(data_mid_68_imag) + $signed(_zz_1170));
  assign _zz_9137 = ($signed(twiddle_factor_table_20_real) * $signed(data_mid_85_real));
  assign _zz_9138 = ($signed(twiddle_factor_table_20_imag) * $signed(data_mid_85_imag));
  assign _zz_9139 = fixTo_586_dout;
  assign _zz_9140 = ($signed(twiddle_factor_table_20_real) * $signed(data_mid_85_imag));
  assign _zz_9141 = ($signed(twiddle_factor_table_20_imag) * $signed(data_mid_85_real));
  assign _zz_9142 = fixTo_587_dout;
  assign _zz_9143 = _zz_9144;
  assign _zz_9144 = ($signed(_zz_9145) >>> _zz_1175);
  assign _zz_9145 = _zz_9146;
  assign _zz_9146 = ($signed(data_mid_69_real) - $signed(_zz_1173));
  assign _zz_9147 = _zz_9148;
  assign _zz_9148 = ($signed(_zz_9149) >>> _zz_1175);
  assign _zz_9149 = _zz_9150;
  assign _zz_9150 = ($signed(data_mid_69_imag) - $signed(_zz_1174));
  assign _zz_9151 = _zz_9152;
  assign _zz_9152 = ($signed(_zz_9153) >>> _zz_1176);
  assign _zz_9153 = _zz_9154;
  assign _zz_9154 = ($signed(data_mid_69_real) + $signed(_zz_1173));
  assign _zz_9155 = _zz_9156;
  assign _zz_9156 = ($signed(_zz_9157) >>> _zz_1176);
  assign _zz_9157 = _zz_9158;
  assign _zz_9158 = ($signed(data_mid_69_imag) + $signed(_zz_1174));
  assign _zz_9159 = ($signed(twiddle_factor_table_21_real) * $signed(data_mid_86_real));
  assign _zz_9160 = ($signed(twiddle_factor_table_21_imag) * $signed(data_mid_86_imag));
  assign _zz_9161 = fixTo_588_dout;
  assign _zz_9162 = ($signed(twiddle_factor_table_21_real) * $signed(data_mid_86_imag));
  assign _zz_9163 = ($signed(twiddle_factor_table_21_imag) * $signed(data_mid_86_real));
  assign _zz_9164 = fixTo_589_dout;
  assign _zz_9165 = _zz_9166;
  assign _zz_9166 = ($signed(_zz_9167) >>> _zz_1179);
  assign _zz_9167 = _zz_9168;
  assign _zz_9168 = ($signed(data_mid_70_real) - $signed(_zz_1177));
  assign _zz_9169 = _zz_9170;
  assign _zz_9170 = ($signed(_zz_9171) >>> _zz_1179);
  assign _zz_9171 = _zz_9172;
  assign _zz_9172 = ($signed(data_mid_70_imag) - $signed(_zz_1178));
  assign _zz_9173 = _zz_9174;
  assign _zz_9174 = ($signed(_zz_9175) >>> _zz_1180);
  assign _zz_9175 = _zz_9176;
  assign _zz_9176 = ($signed(data_mid_70_real) + $signed(_zz_1177));
  assign _zz_9177 = _zz_9178;
  assign _zz_9178 = ($signed(_zz_9179) >>> _zz_1180);
  assign _zz_9179 = _zz_9180;
  assign _zz_9180 = ($signed(data_mid_70_imag) + $signed(_zz_1178));
  assign _zz_9181 = ($signed(twiddle_factor_table_22_real) * $signed(data_mid_87_real));
  assign _zz_9182 = ($signed(twiddle_factor_table_22_imag) * $signed(data_mid_87_imag));
  assign _zz_9183 = fixTo_590_dout;
  assign _zz_9184 = ($signed(twiddle_factor_table_22_real) * $signed(data_mid_87_imag));
  assign _zz_9185 = ($signed(twiddle_factor_table_22_imag) * $signed(data_mid_87_real));
  assign _zz_9186 = fixTo_591_dout;
  assign _zz_9187 = _zz_9188;
  assign _zz_9188 = ($signed(_zz_9189) >>> _zz_1183);
  assign _zz_9189 = _zz_9190;
  assign _zz_9190 = ($signed(data_mid_71_real) - $signed(_zz_1181));
  assign _zz_9191 = _zz_9192;
  assign _zz_9192 = ($signed(_zz_9193) >>> _zz_1183);
  assign _zz_9193 = _zz_9194;
  assign _zz_9194 = ($signed(data_mid_71_imag) - $signed(_zz_1182));
  assign _zz_9195 = _zz_9196;
  assign _zz_9196 = ($signed(_zz_9197) >>> _zz_1184);
  assign _zz_9197 = _zz_9198;
  assign _zz_9198 = ($signed(data_mid_71_real) + $signed(_zz_1181));
  assign _zz_9199 = _zz_9200;
  assign _zz_9200 = ($signed(_zz_9201) >>> _zz_1184);
  assign _zz_9201 = _zz_9202;
  assign _zz_9202 = ($signed(data_mid_71_imag) + $signed(_zz_1182));
  assign _zz_9203 = ($signed(twiddle_factor_table_23_real) * $signed(data_mid_88_real));
  assign _zz_9204 = ($signed(twiddle_factor_table_23_imag) * $signed(data_mid_88_imag));
  assign _zz_9205 = fixTo_592_dout;
  assign _zz_9206 = ($signed(twiddle_factor_table_23_real) * $signed(data_mid_88_imag));
  assign _zz_9207 = ($signed(twiddle_factor_table_23_imag) * $signed(data_mid_88_real));
  assign _zz_9208 = fixTo_593_dout;
  assign _zz_9209 = _zz_9210;
  assign _zz_9210 = ($signed(_zz_9211) >>> _zz_1187);
  assign _zz_9211 = _zz_9212;
  assign _zz_9212 = ($signed(data_mid_72_real) - $signed(_zz_1185));
  assign _zz_9213 = _zz_9214;
  assign _zz_9214 = ($signed(_zz_9215) >>> _zz_1187);
  assign _zz_9215 = _zz_9216;
  assign _zz_9216 = ($signed(data_mid_72_imag) - $signed(_zz_1186));
  assign _zz_9217 = _zz_9218;
  assign _zz_9218 = ($signed(_zz_9219) >>> _zz_1188);
  assign _zz_9219 = _zz_9220;
  assign _zz_9220 = ($signed(data_mid_72_real) + $signed(_zz_1185));
  assign _zz_9221 = _zz_9222;
  assign _zz_9222 = ($signed(_zz_9223) >>> _zz_1188);
  assign _zz_9223 = _zz_9224;
  assign _zz_9224 = ($signed(data_mid_72_imag) + $signed(_zz_1186));
  assign _zz_9225 = ($signed(twiddle_factor_table_24_real) * $signed(data_mid_89_real));
  assign _zz_9226 = ($signed(twiddle_factor_table_24_imag) * $signed(data_mid_89_imag));
  assign _zz_9227 = fixTo_594_dout;
  assign _zz_9228 = ($signed(twiddle_factor_table_24_real) * $signed(data_mid_89_imag));
  assign _zz_9229 = ($signed(twiddle_factor_table_24_imag) * $signed(data_mid_89_real));
  assign _zz_9230 = fixTo_595_dout;
  assign _zz_9231 = _zz_9232;
  assign _zz_9232 = ($signed(_zz_9233) >>> _zz_1191);
  assign _zz_9233 = _zz_9234;
  assign _zz_9234 = ($signed(data_mid_73_real) - $signed(_zz_1189));
  assign _zz_9235 = _zz_9236;
  assign _zz_9236 = ($signed(_zz_9237) >>> _zz_1191);
  assign _zz_9237 = _zz_9238;
  assign _zz_9238 = ($signed(data_mid_73_imag) - $signed(_zz_1190));
  assign _zz_9239 = _zz_9240;
  assign _zz_9240 = ($signed(_zz_9241) >>> _zz_1192);
  assign _zz_9241 = _zz_9242;
  assign _zz_9242 = ($signed(data_mid_73_real) + $signed(_zz_1189));
  assign _zz_9243 = _zz_9244;
  assign _zz_9244 = ($signed(_zz_9245) >>> _zz_1192);
  assign _zz_9245 = _zz_9246;
  assign _zz_9246 = ($signed(data_mid_73_imag) + $signed(_zz_1190));
  assign _zz_9247 = ($signed(twiddle_factor_table_25_real) * $signed(data_mid_90_real));
  assign _zz_9248 = ($signed(twiddle_factor_table_25_imag) * $signed(data_mid_90_imag));
  assign _zz_9249 = fixTo_596_dout;
  assign _zz_9250 = ($signed(twiddle_factor_table_25_real) * $signed(data_mid_90_imag));
  assign _zz_9251 = ($signed(twiddle_factor_table_25_imag) * $signed(data_mid_90_real));
  assign _zz_9252 = fixTo_597_dout;
  assign _zz_9253 = _zz_9254;
  assign _zz_9254 = ($signed(_zz_9255) >>> _zz_1195);
  assign _zz_9255 = _zz_9256;
  assign _zz_9256 = ($signed(data_mid_74_real) - $signed(_zz_1193));
  assign _zz_9257 = _zz_9258;
  assign _zz_9258 = ($signed(_zz_9259) >>> _zz_1195);
  assign _zz_9259 = _zz_9260;
  assign _zz_9260 = ($signed(data_mid_74_imag) - $signed(_zz_1194));
  assign _zz_9261 = _zz_9262;
  assign _zz_9262 = ($signed(_zz_9263) >>> _zz_1196);
  assign _zz_9263 = _zz_9264;
  assign _zz_9264 = ($signed(data_mid_74_real) + $signed(_zz_1193));
  assign _zz_9265 = _zz_9266;
  assign _zz_9266 = ($signed(_zz_9267) >>> _zz_1196);
  assign _zz_9267 = _zz_9268;
  assign _zz_9268 = ($signed(data_mid_74_imag) + $signed(_zz_1194));
  assign _zz_9269 = ($signed(twiddle_factor_table_26_real) * $signed(data_mid_91_real));
  assign _zz_9270 = ($signed(twiddle_factor_table_26_imag) * $signed(data_mid_91_imag));
  assign _zz_9271 = fixTo_598_dout;
  assign _zz_9272 = ($signed(twiddle_factor_table_26_real) * $signed(data_mid_91_imag));
  assign _zz_9273 = ($signed(twiddle_factor_table_26_imag) * $signed(data_mid_91_real));
  assign _zz_9274 = fixTo_599_dout;
  assign _zz_9275 = _zz_9276;
  assign _zz_9276 = ($signed(_zz_9277) >>> _zz_1199);
  assign _zz_9277 = _zz_9278;
  assign _zz_9278 = ($signed(data_mid_75_real) - $signed(_zz_1197));
  assign _zz_9279 = _zz_9280;
  assign _zz_9280 = ($signed(_zz_9281) >>> _zz_1199);
  assign _zz_9281 = _zz_9282;
  assign _zz_9282 = ($signed(data_mid_75_imag) - $signed(_zz_1198));
  assign _zz_9283 = _zz_9284;
  assign _zz_9284 = ($signed(_zz_9285) >>> _zz_1200);
  assign _zz_9285 = _zz_9286;
  assign _zz_9286 = ($signed(data_mid_75_real) + $signed(_zz_1197));
  assign _zz_9287 = _zz_9288;
  assign _zz_9288 = ($signed(_zz_9289) >>> _zz_1200);
  assign _zz_9289 = _zz_9290;
  assign _zz_9290 = ($signed(data_mid_75_imag) + $signed(_zz_1198));
  assign _zz_9291 = ($signed(twiddle_factor_table_27_real) * $signed(data_mid_92_real));
  assign _zz_9292 = ($signed(twiddle_factor_table_27_imag) * $signed(data_mid_92_imag));
  assign _zz_9293 = fixTo_600_dout;
  assign _zz_9294 = ($signed(twiddle_factor_table_27_real) * $signed(data_mid_92_imag));
  assign _zz_9295 = ($signed(twiddle_factor_table_27_imag) * $signed(data_mid_92_real));
  assign _zz_9296 = fixTo_601_dout;
  assign _zz_9297 = _zz_9298;
  assign _zz_9298 = ($signed(_zz_9299) >>> _zz_1203);
  assign _zz_9299 = _zz_9300;
  assign _zz_9300 = ($signed(data_mid_76_real) - $signed(_zz_1201));
  assign _zz_9301 = _zz_9302;
  assign _zz_9302 = ($signed(_zz_9303) >>> _zz_1203);
  assign _zz_9303 = _zz_9304;
  assign _zz_9304 = ($signed(data_mid_76_imag) - $signed(_zz_1202));
  assign _zz_9305 = _zz_9306;
  assign _zz_9306 = ($signed(_zz_9307) >>> _zz_1204);
  assign _zz_9307 = _zz_9308;
  assign _zz_9308 = ($signed(data_mid_76_real) + $signed(_zz_1201));
  assign _zz_9309 = _zz_9310;
  assign _zz_9310 = ($signed(_zz_9311) >>> _zz_1204);
  assign _zz_9311 = _zz_9312;
  assign _zz_9312 = ($signed(data_mid_76_imag) + $signed(_zz_1202));
  assign _zz_9313 = ($signed(twiddle_factor_table_28_real) * $signed(data_mid_93_real));
  assign _zz_9314 = ($signed(twiddle_factor_table_28_imag) * $signed(data_mid_93_imag));
  assign _zz_9315 = fixTo_602_dout;
  assign _zz_9316 = ($signed(twiddle_factor_table_28_real) * $signed(data_mid_93_imag));
  assign _zz_9317 = ($signed(twiddle_factor_table_28_imag) * $signed(data_mid_93_real));
  assign _zz_9318 = fixTo_603_dout;
  assign _zz_9319 = _zz_9320;
  assign _zz_9320 = ($signed(_zz_9321) >>> _zz_1207);
  assign _zz_9321 = _zz_9322;
  assign _zz_9322 = ($signed(data_mid_77_real) - $signed(_zz_1205));
  assign _zz_9323 = _zz_9324;
  assign _zz_9324 = ($signed(_zz_9325) >>> _zz_1207);
  assign _zz_9325 = _zz_9326;
  assign _zz_9326 = ($signed(data_mid_77_imag) - $signed(_zz_1206));
  assign _zz_9327 = _zz_9328;
  assign _zz_9328 = ($signed(_zz_9329) >>> _zz_1208);
  assign _zz_9329 = _zz_9330;
  assign _zz_9330 = ($signed(data_mid_77_real) + $signed(_zz_1205));
  assign _zz_9331 = _zz_9332;
  assign _zz_9332 = ($signed(_zz_9333) >>> _zz_1208);
  assign _zz_9333 = _zz_9334;
  assign _zz_9334 = ($signed(data_mid_77_imag) + $signed(_zz_1206));
  assign _zz_9335 = ($signed(twiddle_factor_table_29_real) * $signed(data_mid_94_real));
  assign _zz_9336 = ($signed(twiddle_factor_table_29_imag) * $signed(data_mid_94_imag));
  assign _zz_9337 = fixTo_604_dout;
  assign _zz_9338 = ($signed(twiddle_factor_table_29_real) * $signed(data_mid_94_imag));
  assign _zz_9339 = ($signed(twiddle_factor_table_29_imag) * $signed(data_mid_94_real));
  assign _zz_9340 = fixTo_605_dout;
  assign _zz_9341 = _zz_9342;
  assign _zz_9342 = ($signed(_zz_9343) >>> _zz_1211);
  assign _zz_9343 = _zz_9344;
  assign _zz_9344 = ($signed(data_mid_78_real) - $signed(_zz_1209));
  assign _zz_9345 = _zz_9346;
  assign _zz_9346 = ($signed(_zz_9347) >>> _zz_1211);
  assign _zz_9347 = _zz_9348;
  assign _zz_9348 = ($signed(data_mid_78_imag) - $signed(_zz_1210));
  assign _zz_9349 = _zz_9350;
  assign _zz_9350 = ($signed(_zz_9351) >>> _zz_1212);
  assign _zz_9351 = _zz_9352;
  assign _zz_9352 = ($signed(data_mid_78_real) + $signed(_zz_1209));
  assign _zz_9353 = _zz_9354;
  assign _zz_9354 = ($signed(_zz_9355) >>> _zz_1212);
  assign _zz_9355 = _zz_9356;
  assign _zz_9356 = ($signed(data_mid_78_imag) + $signed(_zz_1210));
  assign _zz_9357 = ($signed(twiddle_factor_table_30_real) * $signed(data_mid_95_real));
  assign _zz_9358 = ($signed(twiddle_factor_table_30_imag) * $signed(data_mid_95_imag));
  assign _zz_9359 = fixTo_606_dout;
  assign _zz_9360 = ($signed(twiddle_factor_table_30_real) * $signed(data_mid_95_imag));
  assign _zz_9361 = ($signed(twiddle_factor_table_30_imag) * $signed(data_mid_95_real));
  assign _zz_9362 = fixTo_607_dout;
  assign _zz_9363 = _zz_9364;
  assign _zz_9364 = ($signed(_zz_9365) >>> _zz_1215);
  assign _zz_9365 = _zz_9366;
  assign _zz_9366 = ($signed(data_mid_79_real) - $signed(_zz_1213));
  assign _zz_9367 = _zz_9368;
  assign _zz_9368 = ($signed(_zz_9369) >>> _zz_1215);
  assign _zz_9369 = _zz_9370;
  assign _zz_9370 = ($signed(data_mid_79_imag) - $signed(_zz_1214));
  assign _zz_9371 = _zz_9372;
  assign _zz_9372 = ($signed(_zz_9373) >>> _zz_1216);
  assign _zz_9373 = _zz_9374;
  assign _zz_9374 = ($signed(data_mid_79_real) + $signed(_zz_1213));
  assign _zz_9375 = _zz_9376;
  assign _zz_9376 = ($signed(_zz_9377) >>> _zz_1216);
  assign _zz_9377 = _zz_9378;
  assign _zz_9378 = ($signed(data_mid_79_imag) + $signed(_zz_1214));
  assign _zz_9379 = ($signed(twiddle_factor_table_15_real) * $signed(data_mid_112_real));
  assign _zz_9380 = ($signed(twiddle_factor_table_15_imag) * $signed(data_mid_112_imag));
  assign _zz_9381 = fixTo_608_dout;
  assign _zz_9382 = ($signed(twiddle_factor_table_15_real) * $signed(data_mid_112_imag));
  assign _zz_9383 = ($signed(twiddle_factor_table_15_imag) * $signed(data_mid_112_real));
  assign _zz_9384 = fixTo_609_dout;
  assign _zz_9385 = _zz_9386;
  assign _zz_9386 = ($signed(_zz_9387) >>> _zz_1219);
  assign _zz_9387 = _zz_9388;
  assign _zz_9388 = ($signed(data_mid_96_real) - $signed(_zz_1217));
  assign _zz_9389 = _zz_9390;
  assign _zz_9390 = ($signed(_zz_9391) >>> _zz_1219);
  assign _zz_9391 = _zz_9392;
  assign _zz_9392 = ($signed(data_mid_96_imag) - $signed(_zz_1218));
  assign _zz_9393 = _zz_9394;
  assign _zz_9394 = ($signed(_zz_9395) >>> _zz_1220);
  assign _zz_9395 = _zz_9396;
  assign _zz_9396 = ($signed(data_mid_96_real) + $signed(_zz_1217));
  assign _zz_9397 = _zz_9398;
  assign _zz_9398 = ($signed(_zz_9399) >>> _zz_1220);
  assign _zz_9399 = _zz_9400;
  assign _zz_9400 = ($signed(data_mid_96_imag) + $signed(_zz_1218));
  assign _zz_9401 = ($signed(twiddle_factor_table_16_real) * $signed(data_mid_113_real));
  assign _zz_9402 = ($signed(twiddle_factor_table_16_imag) * $signed(data_mid_113_imag));
  assign _zz_9403 = fixTo_610_dout;
  assign _zz_9404 = ($signed(twiddle_factor_table_16_real) * $signed(data_mid_113_imag));
  assign _zz_9405 = ($signed(twiddle_factor_table_16_imag) * $signed(data_mid_113_real));
  assign _zz_9406 = fixTo_611_dout;
  assign _zz_9407 = _zz_9408;
  assign _zz_9408 = ($signed(_zz_9409) >>> _zz_1223);
  assign _zz_9409 = _zz_9410;
  assign _zz_9410 = ($signed(data_mid_97_real) - $signed(_zz_1221));
  assign _zz_9411 = _zz_9412;
  assign _zz_9412 = ($signed(_zz_9413) >>> _zz_1223);
  assign _zz_9413 = _zz_9414;
  assign _zz_9414 = ($signed(data_mid_97_imag) - $signed(_zz_1222));
  assign _zz_9415 = _zz_9416;
  assign _zz_9416 = ($signed(_zz_9417) >>> _zz_1224);
  assign _zz_9417 = _zz_9418;
  assign _zz_9418 = ($signed(data_mid_97_real) + $signed(_zz_1221));
  assign _zz_9419 = _zz_9420;
  assign _zz_9420 = ($signed(_zz_9421) >>> _zz_1224);
  assign _zz_9421 = _zz_9422;
  assign _zz_9422 = ($signed(data_mid_97_imag) + $signed(_zz_1222));
  assign _zz_9423 = ($signed(twiddle_factor_table_17_real) * $signed(data_mid_114_real));
  assign _zz_9424 = ($signed(twiddle_factor_table_17_imag) * $signed(data_mid_114_imag));
  assign _zz_9425 = fixTo_612_dout;
  assign _zz_9426 = ($signed(twiddle_factor_table_17_real) * $signed(data_mid_114_imag));
  assign _zz_9427 = ($signed(twiddle_factor_table_17_imag) * $signed(data_mid_114_real));
  assign _zz_9428 = fixTo_613_dout;
  assign _zz_9429 = _zz_9430;
  assign _zz_9430 = ($signed(_zz_9431) >>> _zz_1227);
  assign _zz_9431 = _zz_9432;
  assign _zz_9432 = ($signed(data_mid_98_real) - $signed(_zz_1225));
  assign _zz_9433 = _zz_9434;
  assign _zz_9434 = ($signed(_zz_9435) >>> _zz_1227);
  assign _zz_9435 = _zz_9436;
  assign _zz_9436 = ($signed(data_mid_98_imag) - $signed(_zz_1226));
  assign _zz_9437 = _zz_9438;
  assign _zz_9438 = ($signed(_zz_9439) >>> _zz_1228);
  assign _zz_9439 = _zz_9440;
  assign _zz_9440 = ($signed(data_mid_98_real) + $signed(_zz_1225));
  assign _zz_9441 = _zz_9442;
  assign _zz_9442 = ($signed(_zz_9443) >>> _zz_1228);
  assign _zz_9443 = _zz_9444;
  assign _zz_9444 = ($signed(data_mid_98_imag) + $signed(_zz_1226));
  assign _zz_9445 = ($signed(twiddle_factor_table_18_real) * $signed(data_mid_115_real));
  assign _zz_9446 = ($signed(twiddle_factor_table_18_imag) * $signed(data_mid_115_imag));
  assign _zz_9447 = fixTo_614_dout;
  assign _zz_9448 = ($signed(twiddle_factor_table_18_real) * $signed(data_mid_115_imag));
  assign _zz_9449 = ($signed(twiddle_factor_table_18_imag) * $signed(data_mid_115_real));
  assign _zz_9450 = fixTo_615_dout;
  assign _zz_9451 = _zz_9452;
  assign _zz_9452 = ($signed(_zz_9453) >>> _zz_1231);
  assign _zz_9453 = _zz_9454;
  assign _zz_9454 = ($signed(data_mid_99_real) - $signed(_zz_1229));
  assign _zz_9455 = _zz_9456;
  assign _zz_9456 = ($signed(_zz_9457) >>> _zz_1231);
  assign _zz_9457 = _zz_9458;
  assign _zz_9458 = ($signed(data_mid_99_imag) - $signed(_zz_1230));
  assign _zz_9459 = _zz_9460;
  assign _zz_9460 = ($signed(_zz_9461) >>> _zz_1232);
  assign _zz_9461 = _zz_9462;
  assign _zz_9462 = ($signed(data_mid_99_real) + $signed(_zz_1229));
  assign _zz_9463 = _zz_9464;
  assign _zz_9464 = ($signed(_zz_9465) >>> _zz_1232);
  assign _zz_9465 = _zz_9466;
  assign _zz_9466 = ($signed(data_mid_99_imag) + $signed(_zz_1230));
  assign _zz_9467 = ($signed(twiddle_factor_table_19_real) * $signed(data_mid_116_real));
  assign _zz_9468 = ($signed(twiddle_factor_table_19_imag) * $signed(data_mid_116_imag));
  assign _zz_9469 = fixTo_616_dout;
  assign _zz_9470 = ($signed(twiddle_factor_table_19_real) * $signed(data_mid_116_imag));
  assign _zz_9471 = ($signed(twiddle_factor_table_19_imag) * $signed(data_mid_116_real));
  assign _zz_9472 = fixTo_617_dout;
  assign _zz_9473 = _zz_9474;
  assign _zz_9474 = ($signed(_zz_9475) >>> _zz_1235);
  assign _zz_9475 = _zz_9476;
  assign _zz_9476 = ($signed(data_mid_100_real) - $signed(_zz_1233));
  assign _zz_9477 = _zz_9478;
  assign _zz_9478 = ($signed(_zz_9479) >>> _zz_1235);
  assign _zz_9479 = _zz_9480;
  assign _zz_9480 = ($signed(data_mid_100_imag) - $signed(_zz_1234));
  assign _zz_9481 = _zz_9482;
  assign _zz_9482 = ($signed(_zz_9483) >>> _zz_1236);
  assign _zz_9483 = _zz_9484;
  assign _zz_9484 = ($signed(data_mid_100_real) + $signed(_zz_1233));
  assign _zz_9485 = _zz_9486;
  assign _zz_9486 = ($signed(_zz_9487) >>> _zz_1236);
  assign _zz_9487 = _zz_9488;
  assign _zz_9488 = ($signed(data_mid_100_imag) + $signed(_zz_1234));
  assign _zz_9489 = ($signed(twiddle_factor_table_20_real) * $signed(data_mid_117_real));
  assign _zz_9490 = ($signed(twiddle_factor_table_20_imag) * $signed(data_mid_117_imag));
  assign _zz_9491 = fixTo_618_dout;
  assign _zz_9492 = ($signed(twiddle_factor_table_20_real) * $signed(data_mid_117_imag));
  assign _zz_9493 = ($signed(twiddle_factor_table_20_imag) * $signed(data_mid_117_real));
  assign _zz_9494 = fixTo_619_dout;
  assign _zz_9495 = _zz_9496;
  assign _zz_9496 = ($signed(_zz_9497) >>> _zz_1239);
  assign _zz_9497 = _zz_9498;
  assign _zz_9498 = ($signed(data_mid_101_real) - $signed(_zz_1237));
  assign _zz_9499 = _zz_9500;
  assign _zz_9500 = ($signed(_zz_9501) >>> _zz_1239);
  assign _zz_9501 = _zz_9502;
  assign _zz_9502 = ($signed(data_mid_101_imag) - $signed(_zz_1238));
  assign _zz_9503 = _zz_9504;
  assign _zz_9504 = ($signed(_zz_9505) >>> _zz_1240);
  assign _zz_9505 = _zz_9506;
  assign _zz_9506 = ($signed(data_mid_101_real) + $signed(_zz_1237));
  assign _zz_9507 = _zz_9508;
  assign _zz_9508 = ($signed(_zz_9509) >>> _zz_1240);
  assign _zz_9509 = _zz_9510;
  assign _zz_9510 = ($signed(data_mid_101_imag) + $signed(_zz_1238));
  assign _zz_9511 = ($signed(twiddle_factor_table_21_real) * $signed(data_mid_118_real));
  assign _zz_9512 = ($signed(twiddle_factor_table_21_imag) * $signed(data_mid_118_imag));
  assign _zz_9513 = fixTo_620_dout;
  assign _zz_9514 = ($signed(twiddle_factor_table_21_real) * $signed(data_mid_118_imag));
  assign _zz_9515 = ($signed(twiddle_factor_table_21_imag) * $signed(data_mid_118_real));
  assign _zz_9516 = fixTo_621_dout;
  assign _zz_9517 = _zz_9518;
  assign _zz_9518 = ($signed(_zz_9519) >>> _zz_1243);
  assign _zz_9519 = _zz_9520;
  assign _zz_9520 = ($signed(data_mid_102_real) - $signed(_zz_1241));
  assign _zz_9521 = _zz_9522;
  assign _zz_9522 = ($signed(_zz_9523) >>> _zz_1243);
  assign _zz_9523 = _zz_9524;
  assign _zz_9524 = ($signed(data_mid_102_imag) - $signed(_zz_1242));
  assign _zz_9525 = _zz_9526;
  assign _zz_9526 = ($signed(_zz_9527) >>> _zz_1244);
  assign _zz_9527 = _zz_9528;
  assign _zz_9528 = ($signed(data_mid_102_real) + $signed(_zz_1241));
  assign _zz_9529 = _zz_9530;
  assign _zz_9530 = ($signed(_zz_9531) >>> _zz_1244);
  assign _zz_9531 = _zz_9532;
  assign _zz_9532 = ($signed(data_mid_102_imag) + $signed(_zz_1242));
  assign _zz_9533 = ($signed(twiddle_factor_table_22_real) * $signed(data_mid_119_real));
  assign _zz_9534 = ($signed(twiddle_factor_table_22_imag) * $signed(data_mid_119_imag));
  assign _zz_9535 = fixTo_622_dout;
  assign _zz_9536 = ($signed(twiddle_factor_table_22_real) * $signed(data_mid_119_imag));
  assign _zz_9537 = ($signed(twiddle_factor_table_22_imag) * $signed(data_mid_119_real));
  assign _zz_9538 = fixTo_623_dout;
  assign _zz_9539 = _zz_9540;
  assign _zz_9540 = ($signed(_zz_9541) >>> _zz_1247);
  assign _zz_9541 = _zz_9542;
  assign _zz_9542 = ($signed(data_mid_103_real) - $signed(_zz_1245));
  assign _zz_9543 = _zz_9544;
  assign _zz_9544 = ($signed(_zz_9545) >>> _zz_1247);
  assign _zz_9545 = _zz_9546;
  assign _zz_9546 = ($signed(data_mid_103_imag) - $signed(_zz_1246));
  assign _zz_9547 = _zz_9548;
  assign _zz_9548 = ($signed(_zz_9549) >>> _zz_1248);
  assign _zz_9549 = _zz_9550;
  assign _zz_9550 = ($signed(data_mid_103_real) + $signed(_zz_1245));
  assign _zz_9551 = _zz_9552;
  assign _zz_9552 = ($signed(_zz_9553) >>> _zz_1248);
  assign _zz_9553 = _zz_9554;
  assign _zz_9554 = ($signed(data_mid_103_imag) + $signed(_zz_1246));
  assign _zz_9555 = ($signed(twiddle_factor_table_23_real) * $signed(data_mid_120_real));
  assign _zz_9556 = ($signed(twiddle_factor_table_23_imag) * $signed(data_mid_120_imag));
  assign _zz_9557 = fixTo_624_dout;
  assign _zz_9558 = ($signed(twiddle_factor_table_23_real) * $signed(data_mid_120_imag));
  assign _zz_9559 = ($signed(twiddle_factor_table_23_imag) * $signed(data_mid_120_real));
  assign _zz_9560 = fixTo_625_dout;
  assign _zz_9561 = _zz_9562;
  assign _zz_9562 = ($signed(_zz_9563) >>> _zz_1251);
  assign _zz_9563 = _zz_9564;
  assign _zz_9564 = ($signed(data_mid_104_real) - $signed(_zz_1249));
  assign _zz_9565 = _zz_9566;
  assign _zz_9566 = ($signed(_zz_9567) >>> _zz_1251);
  assign _zz_9567 = _zz_9568;
  assign _zz_9568 = ($signed(data_mid_104_imag) - $signed(_zz_1250));
  assign _zz_9569 = _zz_9570;
  assign _zz_9570 = ($signed(_zz_9571) >>> _zz_1252);
  assign _zz_9571 = _zz_9572;
  assign _zz_9572 = ($signed(data_mid_104_real) + $signed(_zz_1249));
  assign _zz_9573 = _zz_9574;
  assign _zz_9574 = ($signed(_zz_9575) >>> _zz_1252);
  assign _zz_9575 = _zz_9576;
  assign _zz_9576 = ($signed(data_mid_104_imag) + $signed(_zz_1250));
  assign _zz_9577 = ($signed(twiddle_factor_table_24_real) * $signed(data_mid_121_real));
  assign _zz_9578 = ($signed(twiddle_factor_table_24_imag) * $signed(data_mid_121_imag));
  assign _zz_9579 = fixTo_626_dout;
  assign _zz_9580 = ($signed(twiddle_factor_table_24_real) * $signed(data_mid_121_imag));
  assign _zz_9581 = ($signed(twiddle_factor_table_24_imag) * $signed(data_mid_121_real));
  assign _zz_9582 = fixTo_627_dout;
  assign _zz_9583 = _zz_9584;
  assign _zz_9584 = ($signed(_zz_9585) >>> _zz_1255);
  assign _zz_9585 = _zz_9586;
  assign _zz_9586 = ($signed(data_mid_105_real) - $signed(_zz_1253));
  assign _zz_9587 = _zz_9588;
  assign _zz_9588 = ($signed(_zz_9589) >>> _zz_1255);
  assign _zz_9589 = _zz_9590;
  assign _zz_9590 = ($signed(data_mid_105_imag) - $signed(_zz_1254));
  assign _zz_9591 = _zz_9592;
  assign _zz_9592 = ($signed(_zz_9593) >>> _zz_1256);
  assign _zz_9593 = _zz_9594;
  assign _zz_9594 = ($signed(data_mid_105_real) + $signed(_zz_1253));
  assign _zz_9595 = _zz_9596;
  assign _zz_9596 = ($signed(_zz_9597) >>> _zz_1256);
  assign _zz_9597 = _zz_9598;
  assign _zz_9598 = ($signed(data_mid_105_imag) + $signed(_zz_1254));
  assign _zz_9599 = ($signed(twiddle_factor_table_25_real) * $signed(data_mid_122_real));
  assign _zz_9600 = ($signed(twiddle_factor_table_25_imag) * $signed(data_mid_122_imag));
  assign _zz_9601 = fixTo_628_dout;
  assign _zz_9602 = ($signed(twiddle_factor_table_25_real) * $signed(data_mid_122_imag));
  assign _zz_9603 = ($signed(twiddle_factor_table_25_imag) * $signed(data_mid_122_real));
  assign _zz_9604 = fixTo_629_dout;
  assign _zz_9605 = _zz_9606;
  assign _zz_9606 = ($signed(_zz_9607) >>> _zz_1259);
  assign _zz_9607 = _zz_9608;
  assign _zz_9608 = ($signed(data_mid_106_real) - $signed(_zz_1257));
  assign _zz_9609 = _zz_9610;
  assign _zz_9610 = ($signed(_zz_9611) >>> _zz_1259);
  assign _zz_9611 = _zz_9612;
  assign _zz_9612 = ($signed(data_mid_106_imag) - $signed(_zz_1258));
  assign _zz_9613 = _zz_9614;
  assign _zz_9614 = ($signed(_zz_9615) >>> _zz_1260);
  assign _zz_9615 = _zz_9616;
  assign _zz_9616 = ($signed(data_mid_106_real) + $signed(_zz_1257));
  assign _zz_9617 = _zz_9618;
  assign _zz_9618 = ($signed(_zz_9619) >>> _zz_1260);
  assign _zz_9619 = _zz_9620;
  assign _zz_9620 = ($signed(data_mid_106_imag) + $signed(_zz_1258));
  assign _zz_9621 = ($signed(twiddle_factor_table_26_real) * $signed(data_mid_123_real));
  assign _zz_9622 = ($signed(twiddle_factor_table_26_imag) * $signed(data_mid_123_imag));
  assign _zz_9623 = fixTo_630_dout;
  assign _zz_9624 = ($signed(twiddle_factor_table_26_real) * $signed(data_mid_123_imag));
  assign _zz_9625 = ($signed(twiddle_factor_table_26_imag) * $signed(data_mid_123_real));
  assign _zz_9626 = fixTo_631_dout;
  assign _zz_9627 = _zz_9628;
  assign _zz_9628 = ($signed(_zz_9629) >>> _zz_1263);
  assign _zz_9629 = _zz_9630;
  assign _zz_9630 = ($signed(data_mid_107_real) - $signed(_zz_1261));
  assign _zz_9631 = _zz_9632;
  assign _zz_9632 = ($signed(_zz_9633) >>> _zz_1263);
  assign _zz_9633 = _zz_9634;
  assign _zz_9634 = ($signed(data_mid_107_imag) - $signed(_zz_1262));
  assign _zz_9635 = _zz_9636;
  assign _zz_9636 = ($signed(_zz_9637) >>> _zz_1264);
  assign _zz_9637 = _zz_9638;
  assign _zz_9638 = ($signed(data_mid_107_real) + $signed(_zz_1261));
  assign _zz_9639 = _zz_9640;
  assign _zz_9640 = ($signed(_zz_9641) >>> _zz_1264);
  assign _zz_9641 = _zz_9642;
  assign _zz_9642 = ($signed(data_mid_107_imag) + $signed(_zz_1262));
  assign _zz_9643 = ($signed(twiddle_factor_table_27_real) * $signed(data_mid_124_real));
  assign _zz_9644 = ($signed(twiddle_factor_table_27_imag) * $signed(data_mid_124_imag));
  assign _zz_9645 = fixTo_632_dout;
  assign _zz_9646 = ($signed(twiddle_factor_table_27_real) * $signed(data_mid_124_imag));
  assign _zz_9647 = ($signed(twiddle_factor_table_27_imag) * $signed(data_mid_124_real));
  assign _zz_9648 = fixTo_633_dout;
  assign _zz_9649 = _zz_9650;
  assign _zz_9650 = ($signed(_zz_9651) >>> _zz_1267);
  assign _zz_9651 = _zz_9652;
  assign _zz_9652 = ($signed(data_mid_108_real) - $signed(_zz_1265));
  assign _zz_9653 = _zz_9654;
  assign _zz_9654 = ($signed(_zz_9655) >>> _zz_1267);
  assign _zz_9655 = _zz_9656;
  assign _zz_9656 = ($signed(data_mid_108_imag) - $signed(_zz_1266));
  assign _zz_9657 = _zz_9658;
  assign _zz_9658 = ($signed(_zz_9659) >>> _zz_1268);
  assign _zz_9659 = _zz_9660;
  assign _zz_9660 = ($signed(data_mid_108_real) + $signed(_zz_1265));
  assign _zz_9661 = _zz_9662;
  assign _zz_9662 = ($signed(_zz_9663) >>> _zz_1268);
  assign _zz_9663 = _zz_9664;
  assign _zz_9664 = ($signed(data_mid_108_imag) + $signed(_zz_1266));
  assign _zz_9665 = ($signed(twiddle_factor_table_28_real) * $signed(data_mid_125_real));
  assign _zz_9666 = ($signed(twiddle_factor_table_28_imag) * $signed(data_mid_125_imag));
  assign _zz_9667 = fixTo_634_dout;
  assign _zz_9668 = ($signed(twiddle_factor_table_28_real) * $signed(data_mid_125_imag));
  assign _zz_9669 = ($signed(twiddle_factor_table_28_imag) * $signed(data_mid_125_real));
  assign _zz_9670 = fixTo_635_dout;
  assign _zz_9671 = _zz_9672;
  assign _zz_9672 = ($signed(_zz_9673) >>> _zz_1271);
  assign _zz_9673 = _zz_9674;
  assign _zz_9674 = ($signed(data_mid_109_real) - $signed(_zz_1269));
  assign _zz_9675 = _zz_9676;
  assign _zz_9676 = ($signed(_zz_9677) >>> _zz_1271);
  assign _zz_9677 = _zz_9678;
  assign _zz_9678 = ($signed(data_mid_109_imag) - $signed(_zz_1270));
  assign _zz_9679 = _zz_9680;
  assign _zz_9680 = ($signed(_zz_9681) >>> _zz_1272);
  assign _zz_9681 = _zz_9682;
  assign _zz_9682 = ($signed(data_mid_109_real) + $signed(_zz_1269));
  assign _zz_9683 = _zz_9684;
  assign _zz_9684 = ($signed(_zz_9685) >>> _zz_1272);
  assign _zz_9685 = _zz_9686;
  assign _zz_9686 = ($signed(data_mid_109_imag) + $signed(_zz_1270));
  assign _zz_9687 = ($signed(twiddle_factor_table_29_real) * $signed(data_mid_126_real));
  assign _zz_9688 = ($signed(twiddle_factor_table_29_imag) * $signed(data_mid_126_imag));
  assign _zz_9689 = fixTo_636_dout;
  assign _zz_9690 = ($signed(twiddle_factor_table_29_real) * $signed(data_mid_126_imag));
  assign _zz_9691 = ($signed(twiddle_factor_table_29_imag) * $signed(data_mid_126_real));
  assign _zz_9692 = fixTo_637_dout;
  assign _zz_9693 = _zz_9694;
  assign _zz_9694 = ($signed(_zz_9695) >>> _zz_1275);
  assign _zz_9695 = _zz_9696;
  assign _zz_9696 = ($signed(data_mid_110_real) - $signed(_zz_1273));
  assign _zz_9697 = _zz_9698;
  assign _zz_9698 = ($signed(_zz_9699) >>> _zz_1275);
  assign _zz_9699 = _zz_9700;
  assign _zz_9700 = ($signed(data_mid_110_imag) - $signed(_zz_1274));
  assign _zz_9701 = _zz_9702;
  assign _zz_9702 = ($signed(_zz_9703) >>> _zz_1276);
  assign _zz_9703 = _zz_9704;
  assign _zz_9704 = ($signed(data_mid_110_real) + $signed(_zz_1273));
  assign _zz_9705 = _zz_9706;
  assign _zz_9706 = ($signed(_zz_9707) >>> _zz_1276);
  assign _zz_9707 = _zz_9708;
  assign _zz_9708 = ($signed(data_mid_110_imag) + $signed(_zz_1274));
  assign _zz_9709 = ($signed(twiddle_factor_table_30_real) * $signed(data_mid_127_real));
  assign _zz_9710 = ($signed(twiddle_factor_table_30_imag) * $signed(data_mid_127_imag));
  assign _zz_9711 = fixTo_638_dout;
  assign _zz_9712 = ($signed(twiddle_factor_table_30_real) * $signed(data_mid_127_imag));
  assign _zz_9713 = ($signed(twiddle_factor_table_30_imag) * $signed(data_mid_127_real));
  assign _zz_9714 = fixTo_639_dout;
  assign _zz_9715 = _zz_9716;
  assign _zz_9716 = ($signed(_zz_9717) >>> _zz_1279);
  assign _zz_9717 = _zz_9718;
  assign _zz_9718 = ($signed(data_mid_111_real) - $signed(_zz_1277));
  assign _zz_9719 = _zz_9720;
  assign _zz_9720 = ($signed(_zz_9721) >>> _zz_1279);
  assign _zz_9721 = _zz_9722;
  assign _zz_9722 = ($signed(data_mid_111_imag) - $signed(_zz_1278));
  assign _zz_9723 = _zz_9724;
  assign _zz_9724 = ($signed(_zz_9725) >>> _zz_1280);
  assign _zz_9725 = _zz_9726;
  assign _zz_9726 = ($signed(data_mid_111_real) + $signed(_zz_1277));
  assign _zz_9727 = _zz_9728;
  assign _zz_9728 = ($signed(_zz_9729) >>> _zz_1280);
  assign _zz_9729 = _zz_9730;
  assign _zz_9730 = ($signed(data_mid_111_imag) + $signed(_zz_1278));
  assign _zz_9731 = ($signed(twiddle_factor_table_31_real) * $signed(data_mid_32_real));
  assign _zz_9732 = ($signed(twiddle_factor_table_31_imag) * $signed(data_mid_32_imag));
  assign _zz_9733 = fixTo_640_dout;
  assign _zz_9734 = ($signed(twiddle_factor_table_31_real) * $signed(data_mid_32_imag));
  assign _zz_9735 = ($signed(twiddle_factor_table_31_imag) * $signed(data_mid_32_real));
  assign _zz_9736 = fixTo_641_dout;
  assign _zz_9737 = _zz_9738;
  assign _zz_9738 = ($signed(_zz_9739) >>> _zz_1283);
  assign _zz_9739 = _zz_9740;
  assign _zz_9740 = ($signed(data_mid_0_real) - $signed(_zz_1281));
  assign _zz_9741 = _zz_9742;
  assign _zz_9742 = ($signed(_zz_9743) >>> _zz_1283);
  assign _zz_9743 = _zz_9744;
  assign _zz_9744 = ($signed(data_mid_0_imag) - $signed(_zz_1282));
  assign _zz_9745 = _zz_9746;
  assign _zz_9746 = ($signed(_zz_9747) >>> _zz_1284);
  assign _zz_9747 = _zz_9748;
  assign _zz_9748 = ($signed(data_mid_0_real) + $signed(_zz_1281));
  assign _zz_9749 = _zz_9750;
  assign _zz_9750 = ($signed(_zz_9751) >>> _zz_1284);
  assign _zz_9751 = _zz_9752;
  assign _zz_9752 = ($signed(data_mid_0_imag) + $signed(_zz_1282));
  assign _zz_9753 = ($signed(twiddle_factor_table_32_real) * $signed(data_mid_33_real));
  assign _zz_9754 = ($signed(twiddle_factor_table_32_imag) * $signed(data_mid_33_imag));
  assign _zz_9755 = fixTo_642_dout;
  assign _zz_9756 = ($signed(twiddle_factor_table_32_real) * $signed(data_mid_33_imag));
  assign _zz_9757 = ($signed(twiddle_factor_table_32_imag) * $signed(data_mid_33_real));
  assign _zz_9758 = fixTo_643_dout;
  assign _zz_9759 = _zz_9760;
  assign _zz_9760 = ($signed(_zz_9761) >>> _zz_1287);
  assign _zz_9761 = _zz_9762;
  assign _zz_9762 = ($signed(data_mid_1_real) - $signed(_zz_1285));
  assign _zz_9763 = _zz_9764;
  assign _zz_9764 = ($signed(_zz_9765) >>> _zz_1287);
  assign _zz_9765 = _zz_9766;
  assign _zz_9766 = ($signed(data_mid_1_imag) - $signed(_zz_1286));
  assign _zz_9767 = _zz_9768;
  assign _zz_9768 = ($signed(_zz_9769) >>> _zz_1288);
  assign _zz_9769 = _zz_9770;
  assign _zz_9770 = ($signed(data_mid_1_real) + $signed(_zz_1285));
  assign _zz_9771 = _zz_9772;
  assign _zz_9772 = ($signed(_zz_9773) >>> _zz_1288);
  assign _zz_9773 = _zz_9774;
  assign _zz_9774 = ($signed(data_mid_1_imag) + $signed(_zz_1286));
  assign _zz_9775 = ($signed(twiddle_factor_table_33_real) * $signed(data_mid_34_real));
  assign _zz_9776 = ($signed(twiddle_factor_table_33_imag) * $signed(data_mid_34_imag));
  assign _zz_9777 = fixTo_644_dout;
  assign _zz_9778 = ($signed(twiddle_factor_table_33_real) * $signed(data_mid_34_imag));
  assign _zz_9779 = ($signed(twiddle_factor_table_33_imag) * $signed(data_mid_34_real));
  assign _zz_9780 = fixTo_645_dout;
  assign _zz_9781 = _zz_9782;
  assign _zz_9782 = ($signed(_zz_9783) >>> _zz_1291);
  assign _zz_9783 = _zz_9784;
  assign _zz_9784 = ($signed(data_mid_2_real) - $signed(_zz_1289));
  assign _zz_9785 = _zz_9786;
  assign _zz_9786 = ($signed(_zz_9787) >>> _zz_1291);
  assign _zz_9787 = _zz_9788;
  assign _zz_9788 = ($signed(data_mid_2_imag) - $signed(_zz_1290));
  assign _zz_9789 = _zz_9790;
  assign _zz_9790 = ($signed(_zz_9791) >>> _zz_1292);
  assign _zz_9791 = _zz_9792;
  assign _zz_9792 = ($signed(data_mid_2_real) + $signed(_zz_1289));
  assign _zz_9793 = _zz_9794;
  assign _zz_9794 = ($signed(_zz_9795) >>> _zz_1292);
  assign _zz_9795 = _zz_9796;
  assign _zz_9796 = ($signed(data_mid_2_imag) + $signed(_zz_1290));
  assign _zz_9797 = ($signed(twiddle_factor_table_34_real) * $signed(data_mid_35_real));
  assign _zz_9798 = ($signed(twiddle_factor_table_34_imag) * $signed(data_mid_35_imag));
  assign _zz_9799 = fixTo_646_dout;
  assign _zz_9800 = ($signed(twiddle_factor_table_34_real) * $signed(data_mid_35_imag));
  assign _zz_9801 = ($signed(twiddle_factor_table_34_imag) * $signed(data_mid_35_real));
  assign _zz_9802 = fixTo_647_dout;
  assign _zz_9803 = _zz_9804;
  assign _zz_9804 = ($signed(_zz_9805) >>> _zz_1295);
  assign _zz_9805 = _zz_9806;
  assign _zz_9806 = ($signed(data_mid_3_real) - $signed(_zz_1293));
  assign _zz_9807 = _zz_9808;
  assign _zz_9808 = ($signed(_zz_9809) >>> _zz_1295);
  assign _zz_9809 = _zz_9810;
  assign _zz_9810 = ($signed(data_mid_3_imag) - $signed(_zz_1294));
  assign _zz_9811 = _zz_9812;
  assign _zz_9812 = ($signed(_zz_9813) >>> _zz_1296);
  assign _zz_9813 = _zz_9814;
  assign _zz_9814 = ($signed(data_mid_3_real) + $signed(_zz_1293));
  assign _zz_9815 = _zz_9816;
  assign _zz_9816 = ($signed(_zz_9817) >>> _zz_1296);
  assign _zz_9817 = _zz_9818;
  assign _zz_9818 = ($signed(data_mid_3_imag) + $signed(_zz_1294));
  assign _zz_9819 = ($signed(twiddle_factor_table_35_real) * $signed(data_mid_36_real));
  assign _zz_9820 = ($signed(twiddle_factor_table_35_imag) * $signed(data_mid_36_imag));
  assign _zz_9821 = fixTo_648_dout;
  assign _zz_9822 = ($signed(twiddle_factor_table_35_real) * $signed(data_mid_36_imag));
  assign _zz_9823 = ($signed(twiddle_factor_table_35_imag) * $signed(data_mid_36_real));
  assign _zz_9824 = fixTo_649_dout;
  assign _zz_9825 = _zz_9826;
  assign _zz_9826 = ($signed(_zz_9827) >>> _zz_1299);
  assign _zz_9827 = _zz_9828;
  assign _zz_9828 = ($signed(data_mid_4_real) - $signed(_zz_1297));
  assign _zz_9829 = _zz_9830;
  assign _zz_9830 = ($signed(_zz_9831) >>> _zz_1299);
  assign _zz_9831 = _zz_9832;
  assign _zz_9832 = ($signed(data_mid_4_imag) - $signed(_zz_1298));
  assign _zz_9833 = _zz_9834;
  assign _zz_9834 = ($signed(_zz_9835) >>> _zz_1300);
  assign _zz_9835 = _zz_9836;
  assign _zz_9836 = ($signed(data_mid_4_real) + $signed(_zz_1297));
  assign _zz_9837 = _zz_9838;
  assign _zz_9838 = ($signed(_zz_9839) >>> _zz_1300);
  assign _zz_9839 = _zz_9840;
  assign _zz_9840 = ($signed(data_mid_4_imag) + $signed(_zz_1298));
  assign _zz_9841 = ($signed(twiddle_factor_table_36_real) * $signed(data_mid_37_real));
  assign _zz_9842 = ($signed(twiddle_factor_table_36_imag) * $signed(data_mid_37_imag));
  assign _zz_9843 = fixTo_650_dout;
  assign _zz_9844 = ($signed(twiddle_factor_table_36_real) * $signed(data_mid_37_imag));
  assign _zz_9845 = ($signed(twiddle_factor_table_36_imag) * $signed(data_mid_37_real));
  assign _zz_9846 = fixTo_651_dout;
  assign _zz_9847 = _zz_9848;
  assign _zz_9848 = ($signed(_zz_9849) >>> _zz_1303);
  assign _zz_9849 = _zz_9850;
  assign _zz_9850 = ($signed(data_mid_5_real) - $signed(_zz_1301));
  assign _zz_9851 = _zz_9852;
  assign _zz_9852 = ($signed(_zz_9853) >>> _zz_1303);
  assign _zz_9853 = _zz_9854;
  assign _zz_9854 = ($signed(data_mid_5_imag) - $signed(_zz_1302));
  assign _zz_9855 = _zz_9856;
  assign _zz_9856 = ($signed(_zz_9857) >>> _zz_1304);
  assign _zz_9857 = _zz_9858;
  assign _zz_9858 = ($signed(data_mid_5_real) + $signed(_zz_1301));
  assign _zz_9859 = _zz_9860;
  assign _zz_9860 = ($signed(_zz_9861) >>> _zz_1304);
  assign _zz_9861 = _zz_9862;
  assign _zz_9862 = ($signed(data_mid_5_imag) + $signed(_zz_1302));
  assign _zz_9863 = ($signed(twiddle_factor_table_37_real) * $signed(data_mid_38_real));
  assign _zz_9864 = ($signed(twiddle_factor_table_37_imag) * $signed(data_mid_38_imag));
  assign _zz_9865 = fixTo_652_dout;
  assign _zz_9866 = ($signed(twiddle_factor_table_37_real) * $signed(data_mid_38_imag));
  assign _zz_9867 = ($signed(twiddle_factor_table_37_imag) * $signed(data_mid_38_real));
  assign _zz_9868 = fixTo_653_dout;
  assign _zz_9869 = _zz_9870;
  assign _zz_9870 = ($signed(_zz_9871) >>> _zz_1307);
  assign _zz_9871 = _zz_9872;
  assign _zz_9872 = ($signed(data_mid_6_real) - $signed(_zz_1305));
  assign _zz_9873 = _zz_9874;
  assign _zz_9874 = ($signed(_zz_9875) >>> _zz_1307);
  assign _zz_9875 = _zz_9876;
  assign _zz_9876 = ($signed(data_mid_6_imag) - $signed(_zz_1306));
  assign _zz_9877 = _zz_9878;
  assign _zz_9878 = ($signed(_zz_9879) >>> _zz_1308);
  assign _zz_9879 = _zz_9880;
  assign _zz_9880 = ($signed(data_mid_6_real) + $signed(_zz_1305));
  assign _zz_9881 = _zz_9882;
  assign _zz_9882 = ($signed(_zz_9883) >>> _zz_1308);
  assign _zz_9883 = _zz_9884;
  assign _zz_9884 = ($signed(data_mid_6_imag) + $signed(_zz_1306));
  assign _zz_9885 = ($signed(twiddle_factor_table_38_real) * $signed(data_mid_39_real));
  assign _zz_9886 = ($signed(twiddle_factor_table_38_imag) * $signed(data_mid_39_imag));
  assign _zz_9887 = fixTo_654_dout;
  assign _zz_9888 = ($signed(twiddle_factor_table_38_real) * $signed(data_mid_39_imag));
  assign _zz_9889 = ($signed(twiddle_factor_table_38_imag) * $signed(data_mid_39_real));
  assign _zz_9890 = fixTo_655_dout;
  assign _zz_9891 = _zz_9892;
  assign _zz_9892 = ($signed(_zz_9893) >>> _zz_1311);
  assign _zz_9893 = _zz_9894;
  assign _zz_9894 = ($signed(data_mid_7_real) - $signed(_zz_1309));
  assign _zz_9895 = _zz_9896;
  assign _zz_9896 = ($signed(_zz_9897) >>> _zz_1311);
  assign _zz_9897 = _zz_9898;
  assign _zz_9898 = ($signed(data_mid_7_imag) - $signed(_zz_1310));
  assign _zz_9899 = _zz_9900;
  assign _zz_9900 = ($signed(_zz_9901) >>> _zz_1312);
  assign _zz_9901 = _zz_9902;
  assign _zz_9902 = ($signed(data_mid_7_real) + $signed(_zz_1309));
  assign _zz_9903 = _zz_9904;
  assign _zz_9904 = ($signed(_zz_9905) >>> _zz_1312);
  assign _zz_9905 = _zz_9906;
  assign _zz_9906 = ($signed(data_mid_7_imag) + $signed(_zz_1310));
  assign _zz_9907 = ($signed(twiddle_factor_table_39_real) * $signed(data_mid_40_real));
  assign _zz_9908 = ($signed(twiddle_factor_table_39_imag) * $signed(data_mid_40_imag));
  assign _zz_9909 = fixTo_656_dout;
  assign _zz_9910 = ($signed(twiddle_factor_table_39_real) * $signed(data_mid_40_imag));
  assign _zz_9911 = ($signed(twiddle_factor_table_39_imag) * $signed(data_mid_40_real));
  assign _zz_9912 = fixTo_657_dout;
  assign _zz_9913 = _zz_9914;
  assign _zz_9914 = ($signed(_zz_9915) >>> _zz_1315);
  assign _zz_9915 = _zz_9916;
  assign _zz_9916 = ($signed(data_mid_8_real) - $signed(_zz_1313));
  assign _zz_9917 = _zz_9918;
  assign _zz_9918 = ($signed(_zz_9919) >>> _zz_1315);
  assign _zz_9919 = _zz_9920;
  assign _zz_9920 = ($signed(data_mid_8_imag) - $signed(_zz_1314));
  assign _zz_9921 = _zz_9922;
  assign _zz_9922 = ($signed(_zz_9923) >>> _zz_1316);
  assign _zz_9923 = _zz_9924;
  assign _zz_9924 = ($signed(data_mid_8_real) + $signed(_zz_1313));
  assign _zz_9925 = _zz_9926;
  assign _zz_9926 = ($signed(_zz_9927) >>> _zz_1316);
  assign _zz_9927 = _zz_9928;
  assign _zz_9928 = ($signed(data_mid_8_imag) + $signed(_zz_1314));
  assign _zz_9929 = ($signed(twiddle_factor_table_40_real) * $signed(data_mid_41_real));
  assign _zz_9930 = ($signed(twiddle_factor_table_40_imag) * $signed(data_mid_41_imag));
  assign _zz_9931 = fixTo_658_dout;
  assign _zz_9932 = ($signed(twiddle_factor_table_40_real) * $signed(data_mid_41_imag));
  assign _zz_9933 = ($signed(twiddle_factor_table_40_imag) * $signed(data_mid_41_real));
  assign _zz_9934 = fixTo_659_dout;
  assign _zz_9935 = _zz_9936;
  assign _zz_9936 = ($signed(_zz_9937) >>> _zz_1319);
  assign _zz_9937 = _zz_9938;
  assign _zz_9938 = ($signed(data_mid_9_real) - $signed(_zz_1317));
  assign _zz_9939 = _zz_9940;
  assign _zz_9940 = ($signed(_zz_9941) >>> _zz_1319);
  assign _zz_9941 = _zz_9942;
  assign _zz_9942 = ($signed(data_mid_9_imag) - $signed(_zz_1318));
  assign _zz_9943 = _zz_9944;
  assign _zz_9944 = ($signed(_zz_9945) >>> _zz_1320);
  assign _zz_9945 = _zz_9946;
  assign _zz_9946 = ($signed(data_mid_9_real) + $signed(_zz_1317));
  assign _zz_9947 = _zz_9948;
  assign _zz_9948 = ($signed(_zz_9949) >>> _zz_1320);
  assign _zz_9949 = _zz_9950;
  assign _zz_9950 = ($signed(data_mid_9_imag) + $signed(_zz_1318));
  assign _zz_9951 = ($signed(twiddle_factor_table_41_real) * $signed(data_mid_42_real));
  assign _zz_9952 = ($signed(twiddle_factor_table_41_imag) * $signed(data_mid_42_imag));
  assign _zz_9953 = fixTo_660_dout;
  assign _zz_9954 = ($signed(twiddle_factor_table_41_real) * $signed(data_mid_42_imag));
  assign _zz_9955 = ($signed(twiddle_factor_table_41_imag) * $signed(data_mid_42_real));
  assign _zz_9956 = fixTo_661_dout;
  assign _zz_9957 = _zz_9958;
  assign _zz_9958 = ($signed(_zz_9959) >>> _zz_1323);
  assign _zz_9959 = _zz_9960;
  assign _zz_9960 = ($signed(data_mid_10_real) - $signed(_zz_1321));
  assign _zz_9961 = _zz_9962;
  assign _zz_9962 = ($signed(_zz_9963) >>> _zz_1323);
  assign _zz_9963 = _zz_9964;
  assign _zz_9964 = ($signed(data_mid_10_imag) - $signed(_zz_1322));
  assign _zz_9965 = _zz_9966;
  assign _zz_9966 = ($signed(_zz_9967) >>> _zz_1324);
  assign _zz_9967 = _zz_9968;
  assign _zz_9968 = ($signed(data_mid_10_real) + $signed(_zz_1321));
  assign _zz_9969 = _zz_9970;
  assign _zz_9970 = ($signed(_zz_9971) >>> _zz_1324);
  assign _zz_9971 = _zz_9972;
  assign _zz_9972 = ($signed(data_mid_10_imag) + $signed(_zz_1322));
  assign _zz_9973 = ($signed(twiddle_factor_table_42_real) * $signed(data_mid_43_real));
  assign _zz_9974 = ($signed(twiddle_factor_table_42_imag) * $signed(data_mid_43_imag));
  assign _zz_9975 = fixTo_662_dout;
  assign _zz_9976 = ($signed(twiddle_factor_table_42_real) * $signed(data_mid_43_imag));
  assign _zz_9977 = ($signed(twiddle_factor_table_42_imag) * $signed(data_mid_43_real));
  assign _zz_9978 = fixTo_663_dout;
  assign _zz_9979 = _zz_9980;
  assign _zz_9980 = ($signed(_zz_9981) >>> _zz_1327);
  assign _zz_9981 = _zz_9982;
  assign _zz_9982 = ($signed(data_mid_11_real) - $signed(_zz_1325));
  assign _zz_9983 = _zz_9984;
  assign _zz_9984 = ($signed(_zz_9985) >>> _zz_1327);
  assign _zz_9985 = _zz_9986;
  assign _zz_9986 = ($signed(data_mid_11_imag) - $signed(_zz_1326));
  assign _zz_9987 = _zz_9988;
  assign _zz_9988 = ($signed(_zz_9989) >>> _zz_1328);
  assign _zz_9989 = _zz_9990;
  assign _zz_9990 = ($signed(data_mid_11_real) + $signed(_zz_1325));
  assign _zz_9991 = _zz_9992;
  assign _zz_9992 = ($signed(_zz_9993) >>> _zz_1328);
  assign _zz_9993 = _zz_9994;
  assign _zz_9994 = ($signed(data_mid_11_imag) + $signed(_zz_1326));
  assign _zz_9995 = ($signed(twiddle_factor_table_43_real) * $signed(data_mid_44_real));
  assign _zz_9996 = ($signed(twiddle_factor_table_43_imag) * $signed(data_mid_44_imag));
  assign _zz_9997 = fixTo_664_dout;
  assign _zz_9998 = ($signed(twiddle_factor_table_43_real) * $signed(data_mid_44_imag));
  assign _zz_9999 = ($signed(twiddle_factor_table_43_imag) * $signed(data_mid_44_real));
  assign _zz_10000 = fixTo_665_dout;
  assign _zz_10001 = _zz_10002;
  assign _zz_10002 = ($signed(_zz_10003) >>> _zz_1331);
  assign _zz_10003 = _zz_10004;
  assign _zz_10004 = ($signed(data_mid_12_real) - $signed(_zz_1329));
  assign _zz_10005 = _zz_10006;
  assign _zz_10006 = ($signed(_zz_10007) >>> _zz_1331);
  assign _zz_10007 = _zz_10008;
  assign _zz_10008 = ($signed(data_mid_12_imag) - $signed(_zz_1330));
  assign _zz_10009 = _zz_10010;
  assign _zz_10010 = ($signed(_zz_10011) >>> _zz_1332);
  assign _zz_10011 = _zz_10012;
  assign _zz_10012 = ($signed(data_mid_12_real) + $signed(_zz_1329));
  assign _zz_10013 = _zz_10014;
  assign _zz_10014 = ($signed(_zz_10015) >>> _zz_1332);
  assign _zz_10015 = _zz_10016;
  assign _zz_10016 = ($signed(data_mid_12_imag) + $signed(_zz_1330));
  assign _zz_10017 = ($signed(twiddle_factor_table_44_real) * $signed(data_mid_45_real));
  assign _zz_10018 = ($signed(twiddle_factor_table_44_imag) * $signed(data_mid_45_imag));
  assign _zz_10019 = fixTo_666_dout;
  assign _zz_10020 = ($signed(twiddle_factor_table_44_real) * $signed(data_mid_45_imag));
  assign _zz_10021 = ($signed(twiddle_factor_table_44_imag) * $signed(data_mid_45_real));
  assign _zz_10022 = fixTo_667_dout;
  assign _zz_10023 = _zz_10024;
  assign _zz_10024 = ($signed(_zz_10025) >>> _zz_1335);
  assign _zz_10025 = _zz_10026;
  assign _zz_10026 = ($signed(data_mid_13_real) - $signed(_zz_1333));
  assign _zz_10027 = _zz_10028;
  assign _zz_10028 = ($signed(_zz_10029) >>> _zz_1335);
  assign _zz_10029 = _zz_10030;
  assign _zz_10030 = ($signed(data_mid_13_imag) - $signed(_zz_1334));
  assign _zz_10031 = _zz_10032;
  assign _zz_10032 = ($signed(_zz_10033) >>> _zz_1336);
  assign _zz_10033 = _zz_10034;
  assign _zz_10034 = ($signed(data_mid_13_real) + $signed(_zz_1333));
  assign _zz_10035 = _zz_10036;
  assign _zz_10036 = ($signed(_zz_10037) >>> _zz_1336);
  assign _zz_10037 = _zz_10038;
  assign _zz_10038 = ($signed(data_mid_13_imag) + $signed(_zz_1334));
  assign _zz_10039 = ($signed(twiddle_factor_table_45_real) * $signed(data_mid_46_real));
  assign _zz_10040 = ($signed(twiddle_factor_table_45_imag) * $signed(data_mid_46_imag));
  assign _zz_10041 = fixTo_668_dout;
  assign _zz_10042 = ($signed(twiddle_factor_table_45_real) * $signed(data_mid_46_imag));
  assign _zz_10043 = ($signed(twiddle_factor_table_45_imag) * $signed(data_mid_46_real));
  assign _zz_10044 = fixTo_669_dout;
  assign _zz_10045 = _zz_10046;
  assign _zz_10046 = ($signed(_zz_10047) >>> _zz_1339);
  assign _zz_10047 = _zz_10048;
  assign _zz_10048 = ($signed(data_mid_14_real) - $signed(_zz_1337));
  assign _zz_10049 = _zz_10050;
  assign _zz_10050 = ($signed(_zz_10051) >>> _zz_1339);
  assign _zz_10051 = _zz_10052;
  assign _zz_10052 = ($signed(data_mid_14_imag) - $signed(_zz_1338));
  assign _zz_10053 = _zz_10054;
  assign _zz_10054 = ($signed(_zz_10055) >>> _zz_1340);
  assign _zz_10055 = _zz_10056;
  assign _zz_10056 = ($signed(data_mid_14_real) + $signed(_zz_1337));
  assign _zz_10057 = _zz_10058;
  assign _zz_10058 = ($signed(_zz_10059) >>> _zz_1340);
  assign _zz_10059 = _zz_10060;
  assign _zz_10060 = ($signed(data_mid_14_imag) + $signed(_zz_1338));
  assign _zz_10061 = ($signed(twiddle_factor_table_46_real) * $signed(data_mid_47_real));
  assign _zz_10062 = ($signed(twiddle_factor_table_46_imag) * $signed(data_mid_47_imag));
  assign _zz_10063 = fixTo_670_dout;
  assign _zz_10064 = ($signed(twiddle_factor_table_46_real) * $signed(data_mid_47_imag));
  assign _zz_10065 = ($signed(twiddle_factor_table_46_imag) * $signed(data_mid_47_real));
  assign _zz_10066 = fixTo_671_dout;
  assign _zz_10067 = _zz_10068;
  assign _zz_10068 = ($signed(_zz_10069) >>> _zz_1343);
  assign _zz_10069 = _zz_10070;
  assign _zz_10070 = ($signed(data_mid_15_real) - $signed(_zz_1341));
  assign _zz_10071 = _zz_10072;
  assign _zz_10072 = ($signed(_zz_10073) >>> _zz_1343);
  assign _zz_10073 = _zz_10074;
  assign _zz_10074 = ($signed(data_mid_15_imag) - $signed(_zz_1342));
  assign _zz_10075 = _zz_10076;
  assign _zz_10076 = ($signed(_zz_10077) >>> _zz_1344);
  assign _zz_10077 = _zz_10078;
  assign _zz_10078 = ($signed(data_mid_15_real) + $signed(_zz_1341));
  assign _zz_10079 = _zz_10080;
  assign _zz_10080 = ($signed(_zz_10081) >>> _zz_1344);
  assign _zz_10081 = _zz_10082;
  assign _zz_10082 = ($signed(data_mid_15_imag) + $signed(_zz_1342));
  assign _zz_10083 = ($signed(twiddle_factor_table_47_real) * $signed(data_mid_48_real));
  assign _zz_10084 = ($signed(twiddle_factor_table_47_imag) * $signed(data_mid_48_imag));
  assign _zz_10085 = fixTo_672_dout;
  assign _zz_10086 = ($signed(twiddle_factor_table_47_real) * $signed(data_mid_48_imag));
  assign _zz_10087 = ($signed(twiddle_factor_table_47_imag) * $signed(data_mid_48_real));
  assign _zz_10088 = fixTo_673_dout;
  assign _zz_10089 = _zz_10090;
  assign _zz_10090 = ($signed(_zz_10091) >>> _zz_1347);
  assign _zz_10091 = _zz_10092;
  assign _zz_10092 = ($signed(data_mid_16_real) - $signed(_zz_1345));
  assign _zz_10093 = _zz_10094;
  assign _zz_10094 = ($signed(_zz_10095) >>> _zz_1347);
  assign _zz_10095 = _zz_10096;
  assign _zz_10096 = ($signed(data_mid_16_imag) - $signed(_zz_1346));
  assign _zz_10097 = _zz_10098;
  assign _zz_10098 = ($signed(_zz_10099) >>> _zz_1348);
  assign _zz_10099 = _zz_10100;
  assign _zz_10100 = ($signed(data_mid_16_real) + $signed(_zz_1345));
  assign _zz_10101 = _zz_10102;
  assign _zz_10102 = ($signed(_zz_10103) >>> _zz_1348);
  assign _zz_10103 = _zz_10104;
  assign _zz_10104 = ($signed(data_mid_16_imag) + $signed(_zz_1346));
  assign _zz_10105 = ($signed(twiddle_factor_table_48_real) * $signed(data_mid_49_real));
  assign _zz_10106 = ($signed(twiddle_factor_table_48_imag) * $signed(data_mid_49_imag));
  assign _zz_10107 = fixTo_674_dout;
  assign _zz_10108 = ($signed(twiddle_factor_table_48_real) * $signed(data_mid_49_imag));
  assign _zz_10109 = ($signed(twiddle_factor_table_48_imag) * $signed(data_mid_49_real));
  assign _zz_10110 = fixTo_675_dout;
  assign _zz_10111 = _zz_10112;
  assign _zz_10112 = ($signed(_zz_10113) >>> _zz_1351);
  assign _zz_10113 = _zz_10114;
  assign _zz_10114 = ($signed(data_mid_17_real) - $signed(_zz_1349));
  assign _zz_10115 = _zz_10116;
  assign _zz_10116 = ($signed(_zz_10117) >>> _zz_1351);
  assign _zz_10117 = _zz_10118;
  assign _zz_10118 = ($signed(data_mid_17_imag) - $signed(_zz_1350));
  assign _zz_10119 = _zz_10120;
  assign _zz_10120 = ($signed(_zz_10121) >>> _zz_1352);
  assign _zz_10121 = _zz_10122;
  assign _zz_10122 = ($signed(data_mid_17_real) + $signed(_zz_1349));
  assign _zz_10123 = _zz_10124;
  assign _zz_10124 = ($signed(_zz_10125) >>> _zz_1352);
  assign _zz_10125 = _zz_10126;
  assign _zz_10126 = ($signed(data_mid_17_imag) + $signed(_zz_1350));
  assign _zz_10127 = ($signed(twiddle_factor_table_49_real) * $signed(data_mid_50_real));
  assign _zz_10128 = ($signed(twiddle_factor_table_49_imag) * $signed(data_mid_50_imag));
  assign _zz_10129 = fixTo_676_dout;
  assign _zz_10130 = ($signed(twiddle_factor_table_49_real) * $signed(data_mid_50_imag));
  assign _zz_10131 = ($signed(twiddle_factor_table_49_imag) * $signed(data_mid_50_real));
  assign _zz_10132 = fixTo_677_dout;
  assign _zz_10133 = _zz_10134;
  assign _zz_10134 = ($signed(_zz_10135) >>> _zz_1355);
  assign _zz_10135 = _zz_10136;
  assign _zz_10136 = ($signed(data_mid_18_real) - $signed(_zz_1353));
  assign _zz_10137 = _zz_10138;
  assign _zz_10138 = ($signed(_zz_10139) >>> _zz_1355);
  assign _zz_10139 = _zz_10140;
  assign _zz_10140 = ($signed(data_mid_18_imag) - $signed(_zz_1354));
  assign _zz_10141 = _zz_10142;
  assign _zz_10142 = ($signed(_zz_10143) >>> _zz_1356);
  assign _zz_10143 = _zz_10144;
  assign _zz_10144 = ($signed(data_mid_18_real) + $signed(_zz_1353));
  assign _zz_10145 = _zz_10146;
  assign _zz_10146 = ($signed(_zz_10147) >>> _zz_1356);
  assign _zz_10147 = _zz_10148;
  assign _zz_10148 = ($signed(data_mid_18_imag) + $signed(_zz_1354));
  assign _zz_10149 = ($signed(twiddle_factor_table_50_real) * $signed(data_mid_51_real));
  assign _zz_10150 = ($signed(twiddle_factor_table_50_imag) * $signed(data_mid_51_imag));
  assign _zz_10151 = fixTo_678_dout;
  assign _zz_10152 = ($signed(twiddle_factor_table_50_real) * $signed(data_mid_51_imag));
  assign _zz_10153 = ($signed(twiddle_factor_table_50_imag) * $signed(data_mid_51_real));
  assign _zz_10154 = fixTo_679_dout;
  assign _zz_10155 = _zz_10156;
  assign _zz_10156 = ($signed(_zz_10157) >>> _zz_1359);
  assign _zz_10157 = _zz_10158;
  assign _zz_10158 = ($signed(data_mid_19_real) - $signed(_zz_1357));
  assign _zz_10159 = _zz_10160;
  assign _zz_10160 = ($signed(_zz_10161) >>> _zz_1359);
  assign _zz_10161 = _zz_10162;
  assign _zz_10162 = ($signed(data_mid_19_imag) - $signed(_zz_1358));
  assign _zz_10163 = _zz_10164;
  assign _zz_10164 = ($signed(_zz_10165) >>> _zz_1360);
  assign _zz_10165 = _zz_10166;
  assign _zz_10166 = ($signed(data_mid_19_real) + $signed(_zz_1357));
  assign _zz_10167 = _zz_10168;
  assign _zz_10168 = ($signed(_zz_10169) >>> _zz_1360);
  assign _zz_10169 = _zz_10170;
  assign _zz_10170 = ($signed(data_mid_19_imag) + $signed(_zz_1358));
  assign _zz_10171 = ($signed(twiddle_factor_table_51_real) * $signed(data_mid_52_real));
  assign _zz_10172 = ($signed(twiddle_factor_table_51_imag) * $signed(data_mid_52_imag));
  assign _zz_10173 = fixTo_680_dout;
  assign _zz_10174 = ($signed(twiddle_factor_table_51_real) * $signed(data_mid_52_imag));
  assign _zz_10175 = ($signed(twiddle_factor_table_51_imag) * $signed(data_mid_52_real));
  assign _zz_10176 = fixTo_681_dout;
  assign _zz_10177 = _zz_10178;
  assign _zz_10178 = ($signed(_zz_10179) >>> _zz_1363);
  assign _zz_10179 = _zz_10180;
  assign _zz_10180 = ($signed(data_mid_20_real) - $signed(_zz_1361));
  assign _zz_10181 = _zz_10182;
  assign _zz_10182 = ($signed(_zz_10183) >>> _zz_1363);
  assign _zz_10183 = _zz_10184;
  assign _zz_10184 = ($signed(data_mid_20_imag) - $signed(_zz_1362));
  assign _zz_10185 = _zz_10186;
  assign _zz_10186 = ($signed(_zz_10187) >>> _zz_1364);
  assign _zz_10187 = _zz_10188;
  assign _zz_10188 = ($signed(data_mid_20_real) + $signed(_zz_1361));
  assign _zz_10189 = _zz_10190;
  assign _zz_10190 = ($signed(_zz_10191) >>> _zz_1364);
  assign _zz_10191 = _zz_10192;
  assign _zz_10192 = ($signed(data_mid_20_imag) + $signed(_zz_1362));
  assign _zz_10193 = ($signed(twiddle_factor_table_52_real) * $signed(data_mid_53_real));
  assign _zz_10194 = ($signed(twiddle_factor_table_52_imag) * $signed(data_mid_53_imag));
  assign _zz_10195 = fixTo_682_dout;
  assign _zz_10196 = ($signed(twiddle_factor_table_52_real) * $signed(data_mid_53_imag));
  assign _zz_10197 = ($signed(twiddle_factor_table_52_imag) * $signed(data_mid_53_real));
  assign _zz_10198 = fixTo_683_dout;
  assign _zz_10199 = _zz_10200;
  assign _zz_10200 = ($signed(_zz_10201) >>> _zz_1367);
  assign _zz_10201 = _zz_10202;
  assign _zz_10202 = ($signed(data_mid_21_real) - $signed(_zz_1365));
  assign _zz_10203 = _zz_10204;
  assign _zz_10204 = ($signed(_zz_10205) >>> _zz_1367);
  assign _zz_10205 = _zz_10206;
  assign _zz_10206 = ($signed(data_mid_21_imag) - $signed(_zz_1366));
  assign _zz_10207 = _zz_10208;
  assign _zz_10208 = ($signed(_zz_10209) >>> _zz_1368);
  assign _zz_10209 = _zz_10210;
  assign _zz_10210 = ($signed(data_mid_21_real) + $signed(_zz_1365));
  assign _zz_10211 = _zz_10212;
  assign _zz_10212 = ($signed(_zz_10213) >>> _zz_1368);
  assign _zz_10213 = _zz_10214;
  assign _zz_10214 = ($signed(data_mid_21_imag) + $signed(_zz_1366));
  assign _zz_10215 = ($signed(twiddle_factor_table_53_real) * $signed(data_mid_54_real));
  assign _zz_10216 = ($signed(twiddle_factor_table_53_imag) * $signed(data_mid_54_imag));
  assign _zz_10217 = fixTo_684_dout;
  assign _zz_10218 = ($signed(twiddle_factor_table_53_real) * $signed(data_mid_54_imag));
  assign _zz_10219 = ($signed(twiddle_factor_table_53_imag) * $signed(data_mid_54_real));
  assign _zz_10220 = fixTo_685_dout;
  assign _zz_10221 = _zz_10222;
  assign _zz_10222 = ($signed(_zz_10223) >>> _zz_1371);
  assign _zz_10223 = _zz_10224;
  assign _zz_10224 = ($signed(data_mid_22_real) - $signed(_zz_1369));
  assign _zz_10225 = _zz_10226;
  assign _zz_10226 = ($signed(_zz_10227) >>> _zz_1371);
  assign _zz_10227 = _zz_10228;
  assign _zz_10228 = ($signed(data_mid_22_imag) - $signed(_zz_1370));
  assign _zz_10229 = _zz_10230;
  assign _zz_10230 = ($signed(_zz_10231) >>> _zz_1372);
  assign _zz_10231 = _zz_10232;
  assign _zz_10232 = ($signed(data_mid_22_real) + $signed(_zz_1369));
  assign _zz_10233 = _zz_10234;
  assign _zz_10234 = ($signed(_zz_10235) >>> _zz_1372);
  assign _zz_10235 = _zz_10236;
  assign _zz_10236 = ($signed(data_mid_22_imag) + $signed(_zz_1370));
  assign _zz_10237 = ($signed(twiddle_factor_table_54_real) * $signed(data_mid_55_real));
  assign _zz_10238 = ($signed(twiddle_factor_table_54_imag) * $signed(data_mid_55_imag));
  assign _zz_10239 = fixTo_686_dout;
  assign _zz_10240 = ($signed(twiddle_factor_table_54_real) * $signed(data_mid_55_imag));
  assign _zz_10241 = ($signed(twiddle_factor_table_54_imag) * $signed(data_mid_55_real));
  assign _zz_10242 = fixTo_687_dout;
  assign _zz_10243 = _zz_10244;
  assign _zz_10244 = ($signed(_zz_10245) >>> _zz_1375);
  assign _zz_10245 = _zz_10246;
  assign _zz_10246 = ($signed(data_mid_23_real) - $signed(_zz_1373));
  assign _zz_10247 = _zz_10248;
  assign _zz_10248 = ($signed(_zz_10249) >>> _zz_1375);
  assign _zz_10249 = _zz_10250;
  assign _zz_10250 = ($signed(data_mid_23_imag) - $signed(_zz_1374));
  assign _zz_10251 = _zz_10252;
  assign _zz_10252 = ($signed(_zz_10253) >>> _zz_1376);
  assign _zz_10253 = _zz_10254;
  assign _zz_10254 = ($signed(data_mid_23_real) + $signed(_zz_1373));
  assign _zz_10255 = _zz_10256;
  assign _zz_10256 = ($signed(_zz_10257) >>> _zz_1376);
  assign _zz_10257 = _zz_10258;
  assign _zz_10258 = ($signed(data_mid_23_imag) + $signed(_zz_1374));
  assign _zz_10259 = ($signed(twiddle_factor_table_55_real) * $signed(data_mid_56_real));
  assign _zz_10260 = ($signed(twiddle_factor_table_55_imag) * $signed(data_mid_56_imag));
  assign _zz_10261 = fixTo_688_dout;
  assign _zz_10262 = ($signed(twiddle_factor_table_55_real) * $signed(data_mid_56_imag));
  assign _zz_10263 = ($signed(twiddle_factor_table_55_imag) * $signed(data_mid_56_real));
  assign _zz_10264 = fixTo_689_dout;
  assign _zz_10265 = _zz_10266;
  assign _zz_10266 = ($signed(_zz_10267) >>> _zz_1379);
  assign _zz_10267 = _zz_10268;
  assign _zz_10268 = ($signed(data_mid_24_real) - $signed(_zz_1377));
  assign _zz_10269 = _zz_10270;
  assign _zz_10270 = ($signed(_zz_10271) >>> _zz_1379);
  assign _zz_10271 = _zz_10272;
  assign _zz_10272 = ($signed(data_mid_24_imag) - $signed(_zz_1378));
  assign _zz_10273 = _zz_10274;
  assign _zz_10274 = ($signed(_zz_10275) >>> _zz_1380);
  assign _zz_10275 = _zz_10276;
  assign _zz_10276 = ($signed(data_mid_24_real) + $signed(_zz_1377));
  assign _zz_10277 = _zz_10278;
  assign _zz_10278 = ($signed(_zz_10279) >>> _zz_1380);
  assign _zz_10279 = _zz_10280;
  assign _zz_10280 = ($signed(data_mid_24_imag) + $signed(_zz_1378));
  assign _zz_10281 = ($signed(twiddle_factor_table_56_real) * $signed(data_mid_57_real));
  assign _zz_10282 = ($signed(twiddle_factor_table_56_imag) * $signed(data_mid_57_imag));
  assign _zz_10283 = fixTo_690_dout;
  assign _zz_10284 = ($signed(twiddle_factor_table_56_real) * $signed(data_mid_57_imag));
  assign _zz_10285 = ($signed(twiddle_factor_table_56_imag) * $signed(data_mid_57_real));
  assign _zz_10286 = fixTo_691_dout;
  assign _zz_10287 = _zz_10288;
  assign _zz_10288 = ($signed(_zz_10289) >>> _zz_1383);
  assign _zz_10289 = _zz_10290;
  assign _zz_10290 = ($signed(data_mid_25_real) - $signed(_zz_1381));
  assign _zz_10291 = _zz_10292;
  assign _zz_10292 = ($signed(_zz_10293) >>> _zz_1383);
  assign _zz_10293 = _zz_10294;
  assign _zz_10294 = ($signed(data_mid_25_imag) - $signed(_zz_1382));
  assign _zz_10295 = _zz_10296;
  assign _zz_10296 = ($signed(_zz_10297) >>> _zz_1384);
  assign _zz_10297 = _zz_10298;
  assign _zz_10298 = ($signed(data_mid_25_real) + $signed(_zz_1381));
  assign _zz_10299 = _zz_10300;
  assign _zz_10300 = ($signed(_zz_10301) >>> _zz_1384);
  assign _zz_10301 = _zz_10302;
  assign _zz_10302 = ($signed(data_mid_25_imag) + $signed(_zz_1382));
  assign _zz_10303 = ($signed(twiddle_factor_table_57_real) * $signed(data_mid_58_real));
  assign _zz_10304 = ($signed(twiddle_factor_table_57_imag) * $signed(data_mid_58_imag));
  assign _zz_10305 = fixTo_692_dout;
  assign _zz_10306 = ($signed(twiddle_factor_table_57_real) * $signed(data_mid_58_imag));
  assign _zz_10307 = ($signed(twiddle_factor_table_57_imag) * $signed(data_mid_58_real));
  assign _zz_10308 = fixTo_693_dout;
  assign _zz_10309 = _zz_10310;
  assign _zz_10310 = ($signed(_zz_10311) >>> _zz_1387);
  assign _zz_10311 = _zz_10312;
  assign _zz_10312 = ($signed(data_mid_26_real) - $signed(_zz_1385));
  assign _zz_10313 = _zz_10314;
  assign _zz_10314 = ($signed(_zz_10315) >>> _zz_1387);
  assign _zz_10315 = _zz_10316;
  assign _zz_10316 = ($signed(data_mid_26_imag) - $signed(_zz_1386));
  assign _zz_10317 = _zz_10318;
  assign _zz_10318 = ($signed(_zz_10319) >>> _zz_1388);
  assign _zz_10319 = _zz_10320;
  assign _zz_10320 = ($signed(data_mid_26_real) + $signed(_zz_1385));
  assign _zz_10321 = _zz_10322;
  assign _zz_10322 = ($signed(_zz_10323) >>> _zz_1388);
  assign _zz_10323 = _zz_10324;
  assign _zz_10324 = ($signed(data_mid_26_imag) + $signed(_zz_1386));
  assign _zz_10325 = ($signed(twiddle_factor_table_58_real) * $signed(data_mid_59_real));
  assign _zz_10326 = ($signed(twiddle_factor_table_58_imag) * $signed(data_mid_59_imag));
  assign _zz_10327 = fixTo_694_dout;
  assign _zz_10328 = ($signed(twiddle_factor_table_58_real) * $signed(data_mid_59_imag));
  assign _zz_10329 = ($signed(twiddle_factor_table_58_imag) * $signed(data_mid_59_real));
  assign _zz_10330 = fixTo_695_dout;
  assign _zz_10331 = _zz_10332;
  assign _zz_10332 = ($signed(_zz_10333) >>> _zz_1391);
  assign _zz_10333 = _zz_10334;
  assign _zz_10334 = ($signed(data_mid_27_real) - $signed(_zz_1389));
  assign _zz_10335 = _zz_10336;
  assign _zz_10336 = ($signed(_zz_10337) >>> _zz_1391);
  assign _zz_10337 = _zz_10338;
  assign _zz_10338 = ($signed(data_mid_27_imag) - $signed(_zz_1390));
  assign _zz_10339 = _zz_10340;
  assign _zz_10340 = ($signed(_zz_10341) >>> _zz_1392);
  assign _zz_10341 = _zz_10342;
  assign _zz_10342 = ($signed(data_mid_27_real) + $signed(_zz_1389));
  assign _zz_10343 = _zz_10344;
  assign _zz_10344 = ($signed(_zz_10345) >>> _zz_1392);
  assign _zz_10345 = _zz_10346;
  assign _zz_10346 = ($signed(data_mid_27_imag) + $signed(_zz_1390));
  assign _zz_10347 = ($signed(twiddle_factor_table_59_real) * $signed(data_mid_60_real));
  assign _zz_10348 = ($signed(twiddle_factor_table_59_imag) * $signed(data_mid_60_imag));
  assign _zz_10349 = fixTo_696_dout;
  assign _zz_10350 = ($signed(twiddle_factor_table_59_real) * $signed(data_mid_60_imag));
  assign _zz_10351 = ($signed(twiddle_factor_table_59_imag) * $signed(data_mid_60_real));
  assign _zz_10352 = fixTo_697_dout;
  assign _zz_10353 = _zz_10354;
  assign _zz_10354 = ($signed(_zz_10355) >>> _zz_1395);
  assign _zz_10355 = _zz_10356;
  assign _zz_10356 = ($signed(data_mid_28_real) - $signed(_zz_1393));
  assign _zz_10357 = _zz_10358;
  assign _zz_10358 = ($signed(_zz_10359) >>> _zz_1395);
  assign _zz_10359 = _zz_10360;
  assign _zz_10360 = ($signed(data_mid_28_imag) - $signed(_zz_1394));
  assign _zz_10361 = _zz_10362;
  assign _zz_10362 = ($signed(_zz_10363) >>> _zz_1396);
  assign _zz_10363 = _zz_10364;
  assign _zz_10364 = ($signed(data_mid_28_real) + $signed(_zz_1393));
  assign _zz_10365 = _zz_10366;
  assign _zz_10366 = ($signed(_zz_10367) >>> _zz_1396);
  assign _zz_10367 = _zz_10368;
  assign _zz_10368 = ($signed(data_mid_28_imag) + $signed(_zz_1394));
  assign _zz_10369 = ($signed(twiddle_factor_table_60_real) * $signed(data_mid_61_real));
  assign _zz_10370 = ($signed(twiddle_factor_table_60_imag) * $signed(data_mid_61_imag));
  assign _zz_10371 = fixTo_698_dout;
  assign _zz_10372 = ($signed(twiddle_factor_table_60_real) * $signed(data_mid_61_imag));
  assign _zz_10373 = ($signed(twiddle_factor_table_60_imag) * $signed(data_mid_61_real));
  assign _zz_10374 = fixTo_699_dout;
  assign _zz_10375 = _zz_10376;
  assign _zz_10376 = ($signed(_zz_10377) >>> _zz_1399);
  assign _zz_10377 = _zz_10378;
  assign _zz_10378 = ($signed(data_mid_29_real) - $signed(_zz_1397));
  assign _zz_10379 = _zz_10380;
  assign _zz_10380 = ($signed(_zz_10381) >>> _zz_1399);
  assign _zz_10381 = _zz_10382;
  assign _zz_10382 = ($signed(data_mid_29_imag) - $signed(_zz_1398));
  assign _zz_10383 = _zz_10384;
  assign _zz_10384 = ($signed(_zz_10385) >>> _zz_1400);
  assign _zz_10385 = _zz_10386;
  assign _zz_10386 = ($signed(data_mid_29_real) + $signed(_zz_1397));
  assign _zz_10387 = _zz_10388;
  assign _zz_10388 = ($signed(_zz_10389) >>> _zz_1400);
  assign _zz_10389 = _zz_10390;
  assign _zz_10390 = ($signed(data_mid_29_imag) + $signed(_zz_1398));
  assign _zz_10391 = ($signed(twiddle_factor_table_61_real) * $signed(data_mid_62_real));
  assign _zz_10392 = ($signed(twiddle_factor_table_61_imag) * $signed(data_mid_62_imag));
  assign _zz_10393 = fixTo_700_dout;
  assign _zz_10394 = ($signed(twiddle_factor_table_61_real) * $signed(data_mid_62_imag));
  assign _zz_10395 = ($signed(twiddle_factor_table_61_imag) * $signed(data_mid_62_real));
  assign _zz_10396 = fixTo_701_dout;
  assign _zz_10397 = _zz_10398;
  assign _zz_10398 = ($signed(_zz_10399) >>> _zz_1403);
  assign _zz_10399 = _zz_10400;
  assign _zz_10400 = ($signed(data_mid_30_real) - $signed(_zz_1401));
  assign _zz_10401 = _zz_10402;
  assign _zz_10402 = ($signed(_zz_10403) >>> _zz_1403);
  assign _zz_10403 = _zz_10404;
  assign _zz_10404 = ($signed(data_mid_30_imag) - $signed(_zz_1402));
  assign _zz_10405 = _zz_10406;
  assign _zz_10406 = ($signed(_zz_10407) >>> _zz_1404);
  assign _zz_10407 = _zz_10408;
  assign _zz_10408 = ($signed(data_mid_30_real) + $signed(_zz_1401));
  assign _zz_10409 = _zz_10410;
  assign _zz_10410 = ($signed(_zz_10411) >>> _zz_1404);
  assign _zz_10411 = _zz_10412;
  assign _zz_10412 = ($signed(data_mid_30_imag) + $signed(_zz_1402));
  assign _zz_10413 = ($signed(twiddle_factor_table_62_real) * $signed(data_mid_63_real));
  assign _zz_10414 = ($signed(twiddle_factor_table_62_imag) * $signed(data_mid_63_imag));
  assign _zz_10415 = fixTo_702_dout;
  assign _zz_10416 = ($signed(twiddle_factor_table_62_real) * $signed(data_mid_63_imag));
  assign _zz_10417 = ($signed(twiddle_factor_table_62_imag) * $signed(data_mid_63_real));
  assign _zz_10418 = fixTo_703_dout;
  assign _zz_10419 = _zz_10420;
  assign _zz_10420 = ($signed(_zz_10421) >>> _zz_1407);
  assign _zz_10421 = _zz_10422;
  assign _zz_10422 = ($signed(data_mid_31_real) - $signed(_zz_1405));
  assign _zz_10423 = _zz_10424;
  assign _zz_10424 = ($signed(_zz_10425) >>> _zz_1407);
  assign _zz_10425 = _zz_10426;
  assign _zz_10426 = ($signed(data_mid_31_imag) - $signed(_zz_1406));
  assign _zz_10427 = _zz_10428;
  assign _zz_10428 = ($signed(_zz_10429) >>> _zz_1408);
  assign _zz_10429 = _zz_10430;
  assign _zz_10430 = ($signed(data_mid_31_real) + $signed(_zz_1405));
  assign _zz_10431 = _zz_10432;
  assign _zz_10432 = ($signed(_zz_10433) >>> _zz_1408);
  assign _zz_10433 = _zz_10434;
  assign _zz_10434 = ($signed(data_mid_31_imag) + $signed(_zz_1406));
  assign _zz_10435 = ($signed(twiddle_factor_table_31_real) * $signed(data_mid_96_real));
  assign _zz_10436 = ($signed(twiddle_factor_table_31_imag) * $signed(data_mid_96_imag));
  assign _zz_10437 = fixTo_704_dout;
  assign _zz_10438 = ($signed(twiddle_factor_table_31_real) * $signed(data_mid_96_imag));
  assign _zz_10439 = ($signed(twiddle_factor_table_31_imag) * $signed(data_mid_96_real));
  assign _zz_10440 = fixTo_705_dout;
  assign _zz_10441 = _zz_10442;
  assign _zz_10442 = ($signed(_zz_10443) >>> _zz_1411);
  assign _zz_10443 = _zz_10444;
  assign _zz_10444 = ($signed(data_mid_64_real) - $signed(_zz_1409));
  assign _zz_10445 = _zz_10446;
  assign _zz_10446 = ($signed(_zz_10447) >>> _zz_1411);
  assign _zz_10447 = _zz_10448;
  assign _zz_10448 = ($signed(data_mid_64_imag) - $signed(_zz_1410));
  assign _zz_10449 = _zz_10450;
  assign _zz_10450 = ($signed(_zz_10451) >>> _zz_1412);
  assign _zz_10451 = _zz_10452;
  assign _zz_10452 = ($signed(data_mid_64_real) + $signed(_zz_1409));
  assign _zz_10453 = _zz_10454;
  assign _zz_10454 = ($signed(_zz_10455) >>> _zz_1412);
  assign _zz_10455 = _zz_10456;
  assign _zz_10456 = ($signed(data_mid_64_imag) + $signed(_zz_1410));
  assign _zz_10457 = ($signed(twiddle_factor_table_32_real) * $signed(data_mid_97_real));
  assign _zz_10458 = ($signed(twiddle_factor_table_32_imag) * $signed(data_mid_97_imag));
  assign _zz_10459 = fixTo_706_dout;
  assign _zz_10460 = ($signed(twiddle_factor_table_32_real) * $signed(data_mid_97_imag));
  assign _zz_10461 = ($signed(twiddle_factor_table_32_imag) * $signed(data_mid_97_real));
  assign _zz_10462 = fixTo_707_dout;
  assign _zz_10463 = _zz_10464;
  assign _zz_10464 = ($signed(_zz_10465) >>> _zz_1415);
  assign _zz_10465 = _zz_10466;
  assign _zz_10466 = ($signed(data_mid_65_real) - $signed(_zz_1413));
  assign _zz_10467 = _zz_10468;
  assign _zz_10468 = ($signed(_zz_10469) >>> _zz_1415);
  assign _zz_10469 = _zz_10470;
  assign _zz_10470 = ($signed(data_mid_65_imag) - $signed(_zz_1414));
  assign _zz_10471 = _zz_10472;
  assign _zz_10472 = ($signed(_zz_10473) >>> _zz_1416);
  assign _zz_10473 = _zz_10474;
  assign _zz_10474 = ($signed(data_mid_65_real) + $signed(_zz_1413));
  assign _zz_10475 = _zz_10476;
  assign _zz_10476 = ($signed(_zz_10477) >>> _zz_1416);
  assign _zz_10477 = _zz_10478;
  assign _zz_10478 = ($signed(data_mid_65_imag) + $signed(_zz_1414));
  assign _zz_10479 = ($signed(twiddle_factor_table_33_real) * $signed(data_mid_98_real));
  assign _zz_10480 = ($signed(twiddle_factor_table_33_imag) * $signed(data_mid_98_imag));
  assign _zz_10481 = fixTo_708_dout;
  assign _zz_10482 = ($signed(twiddle_factor_table_33_real) * $signed(data_mid_98_imag));
  assign _zz_10483 = ($signed(twiddle_factor_table_33_imag) * $signed(data_mid_98_real));
  assign _zz_10484 = fixTo_709_dout;
  assign _zz_10485 = _zz_10486;
  assign _zz_10486 = ($signed(_zz_10487) >>> _zz_1419);
  assign _zz_10487 = _zz_10488;
  assign _zz_10488 = ($signed(data_mid_66_real) - $signed(_zz_1417));
  assign _zz_10489 = _zz_10490;
  assign _zz_10490 = ($signed(_zz_10491) >>> _zz_1419);
  assign _zz_10491 = _zz_10492;
  assign _zz_10492 = ($signed(data_mid_66_imag) - $signed(_zz_1418));
  assign _zz_10493 = _zz_10494;
  assign _zz_10494 = ($signed(_zz_10495) >>> _zz_1420);
  assign _zz_10495 = _zz_10496;
  assign _zz_10496 = ($signed(data_mid_66_real) + $signed(_zz_1417));
  assign _zz_10497 = _zz_10498;
  assign _zz_10498 = ($signed(_zz_10499) >>> _zz_1420);
  assign _zz_10499 = _zz_10500;
  assign _zz_10500 = ($signed(data_mid_66_imag) + $signed(_zz_1418));
  assign _zz_10501 = ($signed(twiddle_factor_table_34_real) * $signed(data_mid_99_real));
  assign _zz_10502 = ($signed(twiddle_factor_table_34_imag) * $signed(data_mid_99_imag));
  assign _zz_10503 = fixTo_710_dout;
  assign _zz_10504 = ($signed(twiddle_factor_table_34_real) * $signed(data_mid_99_imag));
  assign _zz_10505 = ($signed(twiddle_factor_table_34_imag) * $signed(data_mid_99_real));
  assign _zz_10506 = fixTo_711_dout;
  assign _zz_10507 = _zz_10508;
  assign _zz_10508 = ($signed(_zz_10509) >>> _zz_1423);
  assign _zz_10509 = _zz_10510;
  assign _zz_10510 = ($signed(data_mid_67_real) - $signed(_zz_1421));
  assign _zz_10511 = _zz_10512;
  assign _zz_10512 = ($signed(_zz_10513) >>> _zz_1423);
  assign _zz_10513 = _zz_10514;
  assign _zz_10514 = ($signed(data_mid_67_imag) - $signed(_zz_1422));
  assign _zz_10515 = _zz_10516;
  assign _zz_10516 = ($signed(_zz_10517) >>> _zz_1424);
  assign _zz_10517 = _zz_10518;
  assign _zz_10518 = ($signed(data_mid_67_real) + $signed(_zz_1421));
  assign _zz_10519 = _zz_10520;
  assign _zz_10520 = ($signed(_zz_10521) >>> _zz_1424);
  assign _zz_10521 = _zz_10522;
  assign _zz_10522 = ($signed(data_mid_67_imag) + $signed(_zz_1422));
  assign _zz_10523 = ($signed(twiddle_factor_table_35_real) * $signed(data_mid_100_real));
  assign _zz_10524 = ($signed(twiddle_factor_table_35_imag) * $signed(data_mid_100_imag));
  assign _zz_10525 = fixTo_712_dout;
  assign _zz_10526 = ($signed(twiddle_factor_table_35_real) * $signed(data_mid_100_imag));
  assign _zz_10527 = ($signed(twiddle_factor_table_35_imag) * $signed(data_mid_100_real));
  assign _zz_10528 = fixTo_713_dout;
  assign _zz_10529 = _zz_10530;
  assign _zz_10530 = ($signed(_zz_10531) >>> _zz_1427);
  assign _zz_10531 = _zz_10532;
  assign _zz_10532 = ($signed(data_mid_68_real) - $signed(_zz_1425));
  assign _zz_10533 = _zz_10534;
  assign _zz_10534 = ($signed(_zz_10535) >>> _zz_1427);
  assign _zz_10535 = _zz_10536;
  assign _zz_10536 = ($signed(data_mid_68_imag) - $signed(_zz_1426));
  assign _zz_10537 = _zz_10538;
  assign _zz_10538 = ($signed(_zz_10539) >>> _zz_1428);
  assign _zz_10539 = _zz_10540;
  assign _zz_10540 = ($signed(data_mid_68_real) + $signed(_zz_1425));
  assign _zz_10541 = _zz_10542;
  assign _zz_10542 = ($signed(_zz_10543) >>> _zz_1428);
  assign _zz_10543 = _zz_10544;
  assign _zz_10544 = ($signed(data_mid_68_imag) + $signed(_zz_1426));
  assign _zz_10545 = ($signed(twiddle_factor_table_36_real) * $signed(data_mid_101_real));
  assign _zz_10546 = ($signed(twiddle_factor_table_36_imag) * $signed(data_mid_101_imag));
  assign _zz_10547 = fixTo_714_dout;
  assign _zz_10548 = ($signed(twiddle_factor_table_36_real) * $signed(data_mid_101_imag));
  assign _zz_10549 = ($signed(twiddle_factor_table_36_imag) * $signed(data_mid_101_real));
  assign _zz_10550 = fixTo_715_dout;
  assign _zz_10551 = _zz_10552;
  assign _zz_10552 = ($signed(_zz_10553) >>> _zz_1431);
  assign _zz_10553 = _zz_10554;
  assign _zz_10554 = ($signed(data_mid_69_real) - $signed(_zz_1429));
  assign _zz_10555 = _zz_10556;
  assign _zz_10556 = ($signed(_zz_10557) >>> _zz_1431);
  assign _zz_10557 = _zz_10558;
  assign _zz_10558 = ($signed(data_mid_69_imag) - $signed(_zz_1430));
  assign _zz_10559 = _zz_10560;
  assign _zz_10560 = ($signed(_zz_10561) >>> _zz_1432);
  assign _zz_10561 = _zz_10562;
  assign _zz_10562 = ($signed(data_mid_69_real) + $signed(_zz_1429));
  assign _zz_10563 = _zz_10564;
  assign _zz_10564 = ($signed(_zz_10565) >>> _zz_1432);
  assign _zz_10565 = _zz_10566;
  assign _zz_10566 = ($signed(data_mid_69_imag) + $signed(_zz_1430));
  assign _zz_10567 = ($signed(twiddle_factor_table_37_real) * $signed(data_mid_102_real));
  assign _zz_10568 = ($signed(twiddle_factor_table_37_imag) * $signed(data_mid_102_imag));
  assign _zz_10569 = fixTo_716_dout;
  assign _zz_10570 = ($signed(twiddle_factor_table_37_real) * $signed(data_mid_102_imag));
  assign _zz_10571 = ($signed(twiddle_factor_table_37_imag) * $signed(data_mid_102_real));
  assign _zz_10572 = fixTo_717_dout;
  assign _zz_10573 = _zz_10574;
  assign _zz_10574 = ($signed(_zz_10575) >>> _zz_1435);
  assign _zz_10575 = _zz_10576;
  assign _zz_10576 = ($signed(data_mid_70_real) - $signed(_zz_1433));
  assign _zz_10577 = _zz_10578;
  assign _zz_10578 = ($signed(_zz_10579) >>> _zz_1435);
  assign _zz_10579 = _zz_10580;
  assign _zz_10580 = ($signed(data_mid_70_imag) - $signed(_zz_1434));
  assign _zz_10581 = _zz_10582;
  assign _zz_10582 = ($signed(_zz_10583) >>> _zz_1436);
  assign _zz_10583 = _zz_10584;
  assign _zz_10584 = ($signed(data_mid_70_real) + $signed(_zz_1433));
  assign _zz_10585 = _zz_10586;
  assign _zz_10586 = ($signed(_zz_10587) >>> _zz_1436);
  assign _zz_10587 = _zz_10588;
  assign _zz_10588 = ($signed(data_mid_70_imag) + $signed(_zz_1434));
  assign _zz_10589 = ($signed(twiddle_factor_table_38_real) * $signed(data_mid_103_real));
  assign _zz_10590 = ($signed(twiddle_factor_table_38_imag) * $signed(data_mid_103_imag));
  assign _zz_10591 = fixTo_718_dout;
  assign _zz_10592 = ($signed(twiddle_factor_table_38_real) * $signed(data_mid_103_imag));
  assign _zz_10593 = ($signed(twiddle_factor_table_38_imag) * $signed(data_mid_103_real));
  assign _zz_10594 = fixTo_719_dout;
  assign _zz_10595 = _zz_10596;
  assign _zz_10596 = ($signed(_zz_10597) >>> _zz_1439);
  assign _zz_10597 = _zz_10598;
  assign _zz_10598 = ($signed(data_mid_71_real) - $signed(_zz_1437));
  assign _zz_10599 = _zz_10600;
  assign _zz_10600 = ($signed(_zz_10601) >>> _zz_1439);
  assign _zz_10601 = _zz_10602;
  assign _zz_10602 = ($signed(data_mid_71_imag) - $signed(_zz_1438));
  assign _zz_10603 = _zz_10604;
  assign _zz_10604 = ($signed(_zz_10605) >>> _zz_1440);
  assign _zz_10605 = _zz_10606;
  assign _zz_10606 = ($signed(data_mid_71_real) + $signed(_zz_1437));
  assign _zz_10607 = _zz_10608;
  assign _zz_10608 = ($signed(_zz_10609) >>> _zz_1440);
  assign _zz_10609 = _zz_10610;
  assign _zz_10610 = ($signed(data_mid_71_imag) + $signed(_zz_1438));
  assign _zz_10611 = ($signed(twiddle_factor_table_39_real) * $signed(data_mid_104_real));
  assign _zz_10612 = ($signed(twiddle_factor_table_39_imag) * $signed(data_mid_104_imag));
  assign _zz_10613 = fixTo_720_dout;
  assign _zz_10614 = ($signed(twiddle_factor_table_39_real) * $signed(data_mid_104_imag));
  assign _zz_10615 = ($signed(twiddle_factor_table_39_imag) * $signed(data_mid_104_real));
  assign _zz_10616 = fixTo_721_dout;
  assign _zz_10617 = _zz_10618;
  assign _zz_10618 = ($signed(_zz_10619) >>> _zz_1443);
  assign _zz_10619 = _zz_10620;
  assign _zz_10620 = ($signed(data_mid_72_real) - $signed(_zz_1441));
  assign _zz_10621 = _zz_10622;
  assign _zz_10622 = ($signed(_zz_10623) >>> _zz_1443);
  assign _zz_10623 = _zz_10624;
  assign _zz_10624 = ($signed(data_mid_72_imag) - $signed(_zz_1442));
  assign _zz_10625 = _zz_10626;
  assign _zz_10626 = ($signed(_zz_10627) >>> _zz_1444);
  assign _zz_10627 = _zz_10628;
  assign _zz_10628 = ($signed(data_mid_72_real) + $signed(_zz_1441));
  assign _zz_10629 = _zz_10630;
  assign _zz_10630 = ($signed(_zz_10631) >>> _zz_1444);
  assign _zz_10631 = _zz_10632;
  assign _zz_10632 = ($signed(data_mid_72_imag) + $signed(_zz_1442));
  assign _zz_10633 = ($signed(twiddle_factor_table_40_real) * $signed(data_mid_105_real));
  assign _zz_10634 = ($signed(twiddle_factor_table_40_imag) * $signed(data_mid_105_imag));
  assign _zz_10635 = fixTo_722_dout;
  assign _zz_10636 = ($signed(twiddle_factor_table_40_real) * $signed(data_mid_105_imag));
  assign _zz_10637 = ($signed(twiddle_factor_table_40_imag) * $signed(data_mid_105_real));
  assign _zz_10638 = fixTo_723_dout;
  assign _zz_10639 = _zz_10640;
  assign _zz_10640 = ($signed(_zz_10641) >>> _zz_1447);
  assign _zz_10641 = _zz_10642;
  assign _zz_10642 = ($signed(data_mid_73_real) - $signed(_zz_1445));
  assign _zz_10643 = _zz_10644;
  assign _zz_10644 = ($signed(_zz_10645) >>> _zz_1447);
  assign _zz_10645 = _zz_10646;
  assign _zz_10646 = ($signed(data_mid_73_imag) - $signed(_zz_1446));
  assign _zz_10647 = _zz_10648;
  assign _zz_10648 = ($signed(_zz_10649) >>> _zz_1448);
  assign _zz_10649 = _zz_10650;
  assign _zz_10650 = ($signed(data_mid_73_real) + $signed(_zz_1445));
  assign _zz_10651 = _zz_10652;
  assign _zz_10652 = ($signed(_zz_10653) >>> _zz_1448);
  assign _zz_10653 = _zz_10654;
  assign _zz_10654 = ($signed(data_mid_73_imag) + $signed(_zz_1446));
  assign _zz_10655 = ($signed(twiddle_factor_table_41_real) * $signed(data_mid_106_real));
  assign _zz_10656 = ($signed(twiddle_factor_table_41_imag) * $signed(data_mid_106_imag));
  assign _zz_10657 = fixTo_724_dout;
  assign _zz_10658 = ($signed(twiddle_factor_table_41_real) * $signed(data_mid_106_imag));
  assign _zz_10659 = ($signed(twiddle_factor_table_41_imag) * $signed(data_mid_106_real));
  assign _zz_10660 = fixTo_725_dout;
  assign _zz_10661 = _zz_10662;
  assign _zz_10662 = ($signed(_zz_10663) >>> _zz_1451);
  assign _zz_10663 = _zz_10664;
  assign _zz_10664 = ($signed(data_mid_74_real) - $signed(_zz_1449));
  assign _zz_10665 = _zz_10666;
  assign _zz_10666 = ($signed(_zz_10667) >>> _zz_1451);
  assign _zz_10667 = _zz_10668;
  assign _zz_10668 = ($signed(data_mid_74_imag) - $signed(_zz_1450));
  assign _zz_10669 = _zz_10670;
  assign _zz_10670 = ($signed(_zz_10671) >>> _zz_1452);
  assign _zz_10671 = _zz_10672;
  assign _zz_10672 = ($signed(data_mid_74_real) + $signed(_zz_1449));
  assign _zz_10673 = _zz_10674;
  assign _zz_10674 = ($signed(_zz_10675) >>> _zz_1452);
  assign _zz_10675 = _zz_10676;
  assign _zz_10676 = ($signed(data_mid_74_imag) + $signed(_zz_1450));
  assign _zz_10677 = ($signed(twiddle_factor_table_42_real) * $signed(data_mid_107_real));
  assign _zz_10678 = ($signed(twiddle_factor_table_42_imag) * $signed(data_mid_107_imag));
  assign _zz_10679 = fixTo_726_dout;
  assign _zz_10680 = ($signed(twiddle_factor_table_42_real) * $signed(data_mid_107_imag));
  assign _zz_10681 = ($signed(twiddle_factor_table_42_imag) * $signed(data_mid_107_real));
  assign _zz_10682 = fixTo_727_dout;
  assign _zz_10683 = _zz_10684;
  assign _zz_10684 = ($signed(_zz_10685) >>> _zz_1455);
  assign _zz_10685 = _zz_10686;
  assign _zz_10686 = ($signed(data_mid_75_real) - $signed(_zz_1453));
  assign _zz_10687 = _zz_10688;
  assign _zz_10688 = ($signed(_zz_10689) >>> _zz_1455);
  assign _zz_10689 = _zz_10690;
  assign _zz_10690 = ($signed(data_mid_75_imag) - $signed(_zz_1454));
  assign _zz_10691 = _zz_10692;
  assign _zz_10692 = ($signed(_zz_10693) >>> _zz_1456);
  assign _zz_10693 = _zz_10694;
  assign _zz_10694 = ($signed(data_mid_75_real) + $signed(_zz_1453));
  assign _zz_10695 = _zz_10696;
  assign _zz_10696 = ($signed(_zz_10697) >>> _zz_1456);
  assign _zz_10697 = _zz_10698;
  assign _zz_10698 = ($signed(data_mid_75_imag) + $signed(_zz_1454));
  assign _zz_10699 = ($signed(twiddle_factor_table_43_real) * $signed(data_mid_108_real));
  assign _zz_10700 = ($signed(twiddle_factor_table_43_imag) * $signed(data_mid_108_imag));
  assign _zz_10701 = fixTo_728_dout;
  assign _zz_10702 = ($signed(twiddle_factor_table_43_real) * $signed(data_mid_108_imag));
  assign _zz_10703 = ($signed(twiddle_factor_table_43_imag) * $signed(data_mid_108_real));
  assign _zz_10704 = fixTo_729_dout;
  assign _zz_10705 = _zz_10706;
  assign _zz_10706 = ($signed(_zz_10707) >>> _zz_1459);
  assign _zz_10707 = _zz_10708;
  assign _zz_10708 = ($signed(data_mid_76_real) - $signed(_zz_1457));
  assign _zz_10709 = _zz_10710;
  assign _zz_10710 = ($signed(_zz_10711) >>> _zz_1459);
  assign _zz_10711 = _zz_10712;
  assign _zz_10712 = ($signed(data_mid_76_imag) - $signed(_zz_1458));
  assign _zz_10713 = _zz_10714;
  assign _zz_10714 = ($signed(_zz_10715) >>> _zz_1460);
  assign _zz_10715 = _zz_10716;
  assign _zz_10716 = ($signed(data_mid_76_real) + $signed(_zz_1457));
  assign _zz_10717 = _zz_10718;
  assign _zz_10718 = ($signed(_zz_10719) >>> _zz_1460);
  assign _zz_10719 = _zz_10720;
  assign _zz_10720 = ($signed(data_mid_76_imag) + $signed(_zz_1458));
  assign _zz_10721 = ($signed(twiddle_factor_table_44_real) * $signed(data_mid_109_real));
  assign _zz_10722 = ($signed(twiddle_factor_table_44_imag) * $signed(data_mid_109_imag));
  assign _zz_10723 = fixTo_730_dout;
  assign _zz_10724 = ($signed(twiddle_factor_table_44_real) * $signed(data_mid_109_imag));
  assign _zz_10725 = ($signed(twiddle_factor_table_44_imag) * $signed(data_mid_109_real));
  assign _zz_10726 = fixTo_731_dout;
  assign _zz_10727 = _zz_10728;
  assign _zz_10728 = ($signed(_zz_10729) >>> _zz_1463);
  assign _zz_10729 = _zz_10730;
  assign _zz_10730 = ($signed(data_mid_77_real) - $signed(_zz_1461));
  assign _zz_10731 = _zz_10732;
  assign _zz_10732 = ($signed(_zz_10733) >>> _zz_1463);
  assign _zz_10733 = _zz_10734;
  assign _zz_10734 = ($signed(data_mid_77_imag) - $signed(_zz_1462));
  assign _zz_10735 = _zz_10736;
  assign _zz_10736 = ($signed(_zz_10737) >>> _zz_1464);
  assign _zz_10737 = _zz_10738;
  assign _zz_10738 = ($signed(data_mid_77_real) + $signed(_zz_1461));
  assign _zz_10739 = _zz_10740;
  assign _zz_10740 = ($signed(_zz_10741) >>> _zz_1464);
  assign _zz_10741 = _zz_10742;
  assign _zz_10742 = ($signed(data_mid_77_imag) + $signed(_zz_1462));
  assign _zz_10743 = ($signed(twiddle_factor_table_45_real) * $signed(data_mid_110_real));
  assign _zz_10744 = ($signed(twiddle_factor_table_45_imag) * $signed(data_mid_110_imag));
  assign _zz_10745 = fixTo_732_dout;
  assign _zz_10746 = ($signed(twiddle_factor_table_45_real) * $signed(data_mid_110_imag));
  assign _zz_10747 = ($signed(twiddle_factor_table_45_imag) * $signed(data_mid_110_real));
  assign _zz_10748 = fixTo_733_dout;
  assign _zz_10749 = _zz_10750;
  assign _zz_10750 = ($signed(_zz_10751) >>> _zz_1467);
  assign _zz_10751 = _zz_10752;
  assign _zz_10752 = ($signed(data_mid_78_real) - $signed(_zz_1465));
  assign _zz_10753 = _zz_10754;
  assign _zz_10754 = ($signed(_zz_10755) >>> _zz_1467);
  assign _zz_10755 = _zz_10756;
  assign _zz_10756 = ($signed(data_mid_78_imag) - $signed(_zz_1466));
  assign _zz_10757 = _zz_10758;
  assign _zz_10758 = ($signed(_zz_10759) >>> _zz_1468);
  assign _zz_10759 = _zz_10760;
  assign _zz_10760 = ($signed(data_mid_78_real) + $signed(_zz_1465));
  assign _zz_10761 = _zz_10762;
  assign _zz_10762 = ($signed(_zz_10763) >>> _zz_1468);
  assign _zz_10763 = _zz_10764;
  assign _zz_10764 = ($signed(data_mid_78_imag) + $signed(_zz_1466));
  assign _zz_10765 = ($signed(twiddle_factor_table_46_real) * $signed(data_mid_111_real));
  assign _zz_10766 = ($signed(twiddle_factor_table_46_imag) * $signed(data_mid_111_imag));
  assign _zz_10767 = fixTo_734_dout;
  assign _zz_10768 = ($signed(twiddle_factor_table_46_real) * $signed(data_mid_111_imag));
  assign _zz_10769 = ($signed(twiddle_factor_table_46_imag) * $signed(data_mid_111_real));
  assign _zz_10770 = fixTo_735_dout;
  assign _zz_10771 = _zz_10772;
  assign _zz_10772 = ($signed(_zz_10773) >>> _zz_1471);
  assign _zz_10773 = _zz_10774;
  assign _zz_10774 = ($signed(data_mid_79_real) - $signed(_zz_1469));
  assign _zz_10775 = _zz_10776;
  assign _zz_10776 = ($signed(_zz_10777) >>> _zz_1471);
  assign _zz_10777 = _zz_10778;
  assign _zz_10778 = ($signed(data_mid_79_imag) - $signed(_zz_1470));
  assign _zz_10779 = _zz_10780;
  assign _zz_10780 = ($signed(_zz_10781) >>> _zz_1472);
  assign _zz_10781 = _zz_10782;
  assign _zz_10782 = ($signed(data_mid_79_real) + $signed(_zz_1469));
  assign _zz_10783 = _zz_10784;
  assign _zz_10784 = ($signed(_zz_10785) >>> _zz_1472);
  assign _zz_10785 = _zz_10786;
  assign _zz_10786 = ($signed(data_mid_79_imag) + $signed(_zz_1470));
  assign _zz_10787 = ($signed(twiddle_factor_table_47_real) * $signed(data_mid_112_real));
  assign _zz_10788 = ($signed(twiddle_factor_table_47_imag) * $signed(data_mid_112_imag));
  assign _zz_10789 = fixTo_736_dout;
  assign _zz_10790 = ($signed(twiddle_factor_table_47_real) * $signed(data_mid_112_imag));
  assign _zz_10791 = ($signed(twiddle_factor_table_47_imag) * $signed(data_mid_112_real));
  assign _zz_10792 = fixTo_737_dout;
  assign _zz_10793 = _zz_10794;
  assign _zz_10794 = ($signed(_zz_10795) >>> _zz_1475);
  assign _zz_10795 = _zz_10796;
  assign _zz_10796 = ($signed(data_mid_80_real) - $signed(_zz_1473));
  assign _zz_10797 = _zz_10798;
  assign _zz_10798 = ($signed(_zz_10799) >>> _zz_1475);
  assign _zz_10799 = _zz_10800;
  assign _zz_10800 = ($signed(data_mid_80_imag) - $signed(_zz_1474));
  assign _zz_10801 = _zz_10802;
  assign _zz_10802 = ($signed(_zz_10803) >>> _zz_1476);
  assign _zz_10803 = _zz_10804;
  assign _zz_10804 = ($signed(data_mid_80_real) + $signed(_zz_1473));
  assign _zz_10805 = _zz_10806;
  assign _zz_10806 = ($signed(_zz_10807) >>> _zz_1476);
  assign _zz_10807 = _zz_10808;
  assign _zz_10808 = ($signed(data_mid_80_imag) + $signed(_zz_1474));
  assign _zz_10809 = ($signed(twiddle_factor_table_48_real) * $signed(data_mid_113_real));
  assign _zz_10810 = ($signed(twiddle_factor_table_48_imag) * $signed(data_mid_113_imag));
  assign _zz_10811 = fixTo_738_dout;
  assign _zz_10812 = ($signed(twiddle_factor_table_48_real) * $signed(data_mid_113_imag));
  assign _zz_10813 = ($signed(twiddle_factor_table_48_imag) * $signed(data_mid_113_real));
  assign _zz_10814 = fixTo_739_dout;
  assign _zz_10815 = _zz_10816;
  assign _zz_10816 = ($signed(_zz_10817) >>> _zz_1479);
  assign _zz_10817 = _zz_10818;
  assign _zz_10818 = ($signed(data_mid_81_real) - $signed(_zz_1477));
  assign _zz_10819 = _zz_10820;
  assign _zz_10820 = ($signed(_zz_10821) >>> _zz_1479);
  assign _zz_10821 = _zz_10822;
  assign _zz_10822 = ($signed(data_mid_81_imag) - $signed(_zz_1478));
  assign _zz_10823 = _zz_10824;
  assign _zz_10824 = ($signed(_zz_10825) >>> _zz_1480);
  assign _zz_10825 = _zz_10826;
  assign _zz_10826 = ($signed(data_mid_81_real) + $signed(_zz_1477));
  assign _zz_10827 = _zz_10828;
  assign _zz_10828 = ($signed(_zz_10829) >>> _zz_1480);
  assign _zz_10829 = _zz_10830;
  assign _zz_10830 = ($signed(data_mid_81_imag) + $signed(_zz_1478));
  assign _zz_10831 = ($signed(twiddle_factor_table_49_real) * $signed(data_mid_114_real));
  assign _zz_10832 = ($signed(twiddle_factor_table_49_imag) * $signed(data_mid_114_imag));
  assign _zz_10833 = fixTo_740_dout;
  assign _zz_10834 = ($signed(twiddle_factor_table_49_real) * $signed(data_mid_114_imag));
  assign _zz_10835 = ($signed(twiddle_factor_table_49_imag) * $signed(data_mid_114_real));
  assign _zz_10836 = fixTo_741_dout;
  assign _zz_10837 = _zz_10838;
  assign _zz_10838 = ($signed(_zz_10839) >>> _zz_1483);
  assign _zz_10839 = _zz_10840;
  assign _zz_10840 = ($signed(data_mid_82_real) - $signed(_zz_1481));
  assign _zz_10841 = _zz_10842;
  assign _zz_10842 = ($signed(_zz_10843) >>> _zz_1483);
  assign _zz_10843 = _zz_10844;
  assign _zz_10844 = ($signed(data_mid_82_imag) - $signed(_zz_1482));
  assign _zz_10845 = _zz_10846;
  assign _zz_10846 = ($signed(_zz_10847) >>> _zz_1484);
  assign _zz_10847 = _zz_10848;
  assign _zz_10848 = ($signed(data_mid_82_real) + $signed(_zz_1481));
  assign _zz_10849 = _zz_10850;
  assign _zz_10850 = ($signed(_zz_10851) >>> _zz_1484);
  assign _zz_10851 = _zz_10852;
  assign _zz_10852 = ($signed(data_mid_82_imag) + $signed(_zz_1482));
  assign _zz_10853 = ($signed(twiddle_factor_table_50_real) * $signed(data_mid_115_real));
  assign _zz_10854 = ($signed(twiddle_factor_table_50_imag) * $signed(data_mid_115_imag));
  assign _zz_10855 = fixTo_742_dout;
  assign _zz_10856 = ($signed(twiddle_factor_table_50_real) * $signed(data_mid_115_imag));
  assign _zz_10857 = ($signed(twiddle_factor_table_50_imag) * $signed(data_mid_115_real));
  assign _zz_10858 = fixTo_743_dout;
  assign _zz_10859 = _zz_10860;
  assign _zz_10860 = ($signed(_zz_10861) >>> _zz_1487);
  assign _zz_10861 = _zz_10862;
  assign _zz_10862 = ($signed(data_mid_83_real) - $signed(_zz_1485));
  assign _zz_10863 = _zz_10864;
  assign _zz_10864 = ($signed(_zz_10865) >>> _zz_1487);
  assign _zz_10865 = _zz_10866;
  assign _zz_10866 = ($signed(data_mid_83_imag) - $signed(_zz_1486));
  assign _zz_10867 = _zz_10868;
  assign _zz_10868 = ($signed(_zz_10869) >>> _zz_1488);
  assign _zz_10869 = _zz_10870;
  assign _zz_10870 = ($signed(data_mid_83_real) + $signed(_zz_1485));
  assign _zz_10871 = _zz_10872;
  assign _zz_10872 = ($signed(_zz_10873) >>> _zz_1488);
  assign _zz_10873 = _zz_10874;
  assign _zz_10874 = ($signed(data_mid_83_imag) + $signed(_zz_1486));
  assign _zz_10875 = ($signed(twiddle_factor_table_51_real) * $signed(data_mid_116_real));
  assign _zz_10876 = ($signed(twiddle_factor_table_51_imag) * $signed(data_mid_116_imag));
  assign _zz_10877 = fixTo_744_dout;
  assign _zz_10878 = ($signed(twiddle_factor_table_51_real) * $signed(data_mid_116_imag));
  assign _zz_10879 = ($signed(twiddle_factor_table_51_imag) * $signed(data_mid_116_real));
  assign _zz_10880 = fixTo_745_dout;
  assign _zz_10881 = _zz_10882;
  assign _zz_10882 = ($signed(_zz_10883) >>> _zz_1491);
  assign _zz_10883 = _zz_10884;
  assign _zz_10884 = ($signed(data_mid_84_real) - $signed(_zz_1489));
  assign _zz_10885 = _zz_10886;
  assign _zz_10886 = ($signed(_zz_10887) >>> _zz_1491);
  assign _zz_10887 = _zz_10888;
  assign _zz_10888 = ($signed(data_mid_84_imag) - $signed(_zz_1490));
  assign _zz_10889 = _zz_10890;
  assign _zz_10890 = ($signed(_zz_10891) >>> _zz_1492);
  assign _zz_10891 = _zz_10892;
  assign _zz_10892 = ($signed(data_mid_84_real) + $signed(_zz_1489));
  assign _zz_10893 = _zz_10894;
  assign _zz_10894 = ($signed(_zz_10895) >>> _zz_1492);
  assign _zz_10895 = _zz_10896;
  assign _zz_10896 = ($signed(data_mid_84_imag) + $signed(_zz_1490));
  assign _zz_10897 = ($signed(twiddle_factor_table_52_real) * $signed(data_mid_117_real));
  assign _zz_10898 = ($signed(twiddle_factor_table_52_imag) * $signed(data_mid_117_imag));
  assign _zz_10899 = fixTo_746_dout;
  assign _zz_10900 = ($signed(twiddle_factor_table_52_real) * $signed(data_mid_117_imag));
  assign _zz_10901 = ($signed(twiddle_factor_table_52_imag) * $signed(data_mid_117_real));
  assign _zz_10902 = fixTo_747_dout;
  assign _zz_10903 = _zz_10904;
  assign _zz_10904 = ($signed(_zz_10905) >>> _zz_1495);
  assign _zz_10905 = _zz_10906;
  assign _zz_10906 = ($signed(data_mid_85_real) - $signed(_zz_1493));
  assign _zz_10907 = _zz_10908;
  assign _zz_10908 = ($signed(_zz_10909) >>> _zz_1495);
  assign _zz_10909 = _zz_10910;
  assign _zz_10910 = ($signed(data_mid_85_imag) - $signed(_zz_1494));
  assign _zz_10911 = _zz_10912;
  assign _zz_10912 = ($signed(_zz_10913) >>> _zz_1496);
  assign _zz_10913 = _zz_10914;
  assign _zz_10914 = ($signed(data_mid_85_real) + $signed(_zz_1493));
  assign _zz_10915 = _zz_10916;
  assign _zz_10916 = ($signed(_zz_10917) >>> _zz_1496);
  assign _zz_10917 = _zz_10918;
  assign _zz_10918 = ($signed(data_mid_85_imag) + $signed(_zz_1494));
  assign _zz_10919 = ($signed(twiddle_factor_table_53_real) * $signed(data_mid_118_real));
  assign _zz_10920 = ($signed(twiddle_factor_table_53_imag) * $signed(data_mid_118_imag));
  assign _zz_10921 = fixTo_748_dout;
  assign _zz_10922 = ($signed(twiddle_factor_table_53_real) * $signed(data_mid_118_imag));
  assign _zz_10923 = ($signed(twiddle_factor_table_53_imag) * $signed(data_mid_118_real));
  assign _zz_10924 = fixTo_749_dout;
  assign _zz_10925 = _zz_10926;
  assign _zz_10926 = ($signed(_zz_10927) >>> _zz_1499);
  assign _zz_10927 = _zz_10928;
  assign _zz_10928 = ($signed(data_mid_86_real) - $signed(_zz_1497));
  assign _zz_10929 = _zz_10930;
  assign _zz_10930 = ($signed(_zz_10931) >>> _zz_1499);
  assign _zz_10931 = _zz_10932;
  assign _zz_10932 = ($signed(data_mid_86_imag) - $signed(_zz_1498));
  assign _zz_10933 = _zz_10934;
  assign _zz_10934 = ($signed(_zz_10935) >>> _zz_1500);
  assign _zz_10935 = _zz_10936;
  assign _zz_10936 = ($signed(data_mid_86_real) + $signed(_zz_1497));
  assign _zz_10937 = _zz_10938;
  assign _zz_10938 = ($signed(_zz_10939) >>> _zz_1500);
  assign _zz_10939 = _zz_10940;
  assign _zz_10940 = ($signed(data_mid_86_imag) + $signed(_zz_1498));
  assign _zz_10941 = ($signed(twiddle_factor_table_54_real) * $signed(data_mid_119_real));
  assign _zz_10942 = ($signed(twiddle_factor_table_54_imag) * $signed(data_mid_119_imag));
  assign _zz_10943 = fixTo_750_dout;
  assign _zz_10944 = ($signed(twiddle_factor_table_54_real) * $signed(data_mid_119_imag));
  assign _zz_10945 = ($signed(twiddle_factor_table_54_imag) * $signed(data_mid_119_real));
  assign _zz_10946 = fixTo_751_dout;
  assign _zz_10947 = _zz_10948;
  assign _zz_10948 = ($signed(_zz_10949) >>> _zz_1503);
  assign _zz_10949 = _zz_10950;
  assign _zz_10950 = ($signed(data_mid_87_real) - $signed(_zz_1501));
  assign _zz_10951 = _zz_10952;
  assign _zz_10952 = ($signed(_zz_10953) >>> _zz_1503);
  assign _zz_10953 = _zz_10954;
  assign _zz_10954 = ($signed(data_mid_87_imag) - $signed(_zz_1502));
  assign _zz_10955 = _zz_10956;
  assign _zz_10956 = ($signed(_zz_10957) >>> _zz_1504);
  assign _zz_10957 = _zz_10958;
  assign _zz_10958 = ($signed(data_mid_87_real) + $signed(_zz_1501));
  assign _zz_10959 = _zz_10960;
  assign _zz_10960 = ($signed(_zz_10961) >>> _zz_1504);
  assign _zz_10961 = _zz_10962;
  assign _zz_10962 = ($signed(data_mid_87_imag) + $signed(_zz_1502));
  assign _zz_10963 = ($signed(twiddle_factor_table_55_real) * $signed(data_mid_120_real));
  assign _zz_10964 = ($signed(twiddle_factor_table_55_imag) * $signed(data_mid_120_imag));
  assign _zz_10965 = fixTo_752_dout;
  assign _zz_10966 = ($signed(twiddle_factor_table_55_real) * $signed(data_mid_120_imag));
  assign _zz_10967 = ($signed(twiddle_factor_table_55_imag) * $signed(data_mid_120_real));
  assign _zz_10968 = fixTo_753_dout;
  assign _zz_10969 = _zz_10970;
  assign _zz_10970 = ($signed(_zz_10971) >>> _zz_1507);
  assign _zz_10971 = _zz_10972;
  assign _zz_10972 = ($signed(data_mid_88_real) - $signed(_zz_1505));
  assign _zz_10973 = _zz_10974;
  assign _zz_10974 = ($signed(_zz_10975) >>> _zz_1507);
  assign _zz_10975 = _zz_10976;
  assign _zz_10976 = ($signed(data_mid_88_imag) - $signed(_zz_1506));
  assign _zz_10977 = _zz_10978;
  assign _zz_10978 = ($signed(_zz_10979) >>> _zz_1508);
  assign _zz_10979 = _zz_10980;
  assign _zz_10980 = ($signed(data_mid_88_real) + $signed(_zz_1505));
  assign _zz_10981 = _zz_10982;
  assign _zz_10982 = ($signed(_zz_10983) >>> _zz_1508);
  assign _zz_10983 = _zz_10984;
  assign _zz_10984 = ($signed(data_mid_88_imag) + $signed(_zz_1506));
  assign _zz_10985 = ($signed(twiddle_factor_table_56_real) * $signed(data_mid_121_real));
  assign _zz_10986 = ($signed(twiddle_factor_table_56_imag) * $signed(data_mid_121_imag));
  assign _zz_10987 = fixTo_754_dout;
  assign _zz_10988 = ($signed(twiddle_factor_table_56_real) * $signed(data_mid_121_imag));
  assign _zz_10989 = ($signed(twiddle_factor_table_56_imag) * $signed(data_mid_121_real));
  assign _zz_10990 = fixTo_755_dout;
  assign _zz_10991 = _zz_10992;
  assign _zz_10992 = ($signed(_zz_10993) >>> _zz_1511);
  assign _zz_10993 = _zz_10994;
  assign _zz_10994 = ($signed(data_mid_89_real) - $signed(_zz_1509));
  assign _zz_10995 = _zz_10996;
  assign _zz_10996 = ($signed(_zz_10997) >>> _zz_1511);
  assign _zz_10997 = _zz_10998;
  assign _zz_10998 = ($signed(data_mid_89_imag) - $signed(_zz_1510));
  assign _zz_10999 = _zz_11000;
  assign _zz_11000 = ($signed(_zz_11001) >>> _zz_1512);
  assign _zz_11001 = _zz_11002;
  assign _zz_11002 = ($signed(data_mid_89_real) + $signed(_zz_1509));
  assign _zz_11003 = _zz_11004;
  assign _zz_11004 = ($signed(_zz_11005) >>> _zz_1512);
  assign _zz_11005 = _zz_11006;
  assign _zz_11006 = ($signed(data_mid_89_imag) + $signed(_zz_1510));
  assign _zz_11007 = ($signed(twiddle_factor_table_57_real) * $signed(data_mid_122_real));
  assign _zz_11008 = ($signed(twiddle_factor_table_57_imag) * $signed(data_mid_122_imag));
  assign _zz_11009 = fixTo_756_dout;
  assign _zz_11010 = ($signed(twiddle_factor_table_57_real) * $signed(data_mid_122_imag));
  assign _zz_11011 = ($signed(twiddle_factor_table_57_imag) * $signed(data_mid_122_real));
  assign _zz_11012 = fixTo_757_dout;
  assign _zz_11013 = _zz_11014;
  assign _zz_11014 = ($signed(_zz_11015) >>> _zz_1515);
  assign _zz_11015 = _zz_11016;
  assign _zz_11016 = ($signed(data_mid_90_real) - $signed(_zz_1513));
  assign _zz_11017 = _zz_11018;
  assign _zz_11018 = ($signed(_zz_11019) >>> _zz_1515);
  assign _zz_11019 = _zz_11020;
  assign _zz_11020 = ($signed(data_mid_90_imag) - $signed(_zz_1514));
  assign _zz_11021 = _zz_11022;
  assign _zz_11022 = ($signed(_zz_11023) >>> _zz_1516);
  assign _zz_11023 = _zz_11024;
  assign _zz_11024 = ($signed(data_mid_90_real) + $signed(_zz_1513));
  assign _zz_11025 = _zz_11026;
  assign _zz_11026 = ($signed(_zz_11027) >>> _zz_1516);
  assign _zz_11027 = _zz_11028;
  assign _zz_11028 = ($signed(data_mid_90_imag) + $signed(_zz_1514));
  assign _zz_11029 = ($signed(twiddle_factor_table_58_real) * $signed(data_mid_123_real));
  assign _zz_11030 = ($signed(twiddle_factor_table_58_imag) * $signed(data_mid_123_imag));
  assign _zz_11031 = fixTo_758_dout;
  assign _zz_11032 = ($signed(twiddle_factor_table_58_real) * $signed(data_mid_123_imag));
  assign _zz_11033 = ($signed(twiddle_factor_table_58_imag) * $signed(data_mid_123_real));
  assign _zz_11034 = fixTo_759_dout;
  assign _zz_11035 = _zz_11036;
  assign _zz_11036 = ($signed(_zz_11037) >>> _zz_1519);
  assign _zz_11037 = _zz_11038;
  assign _zz_11038 = ($signed(data_mid_91_real) - $signed(_zz_1517));
  assign _zz_11039 = _zz_11040;
  assign _zz_11040 = ($signed(_zz_11041) >>> _zz_1519);
  assign _zz_11041 = _zz_11042;
  assign _zz_11042 = ($signed(data_mid_91_imag) - $signed(_zz_1518));
  assign _zz_11043 = _zz_11044;
  assign _zz_11044 = ($signed(_zz_11045) >>> _zz_1520);
  assign _zz_11045 = _zz_11046;
  assign _zz_11046 = ($signed(data_mid_91_real) + $signed(_zz_1517));
  assign _zz_11047 = _zz_11048;
  assign _zz_11048 = ($signed(_zz_11049) >>> _zz_1520);
  assign _zz_11049 = _zz_11050;
  assign _zz_11050 = ($signed(data_mid_91_imag) + $signed(_zz_1518));
  assign _zz_11051 = ($signed(twiddle_factor_table_59_real) * $signed(data_mid_124_real));
  assign _zz_11052 = ($signed(twiddle_factor_table_59_imag) * $signed(data_mid_124_imag));
  assign _zz_11053 = fixTo_760_dout;
  assign _zz_11054 = ($signed(twiddle_factor_table_59_real) * $signed(data_mid_124_imag));
  assign _zz_11055 = ($signed(twiddle_factor_table_59_imag) * $signed(data_mid_124_real));
  assign _zz_11056 = fixTo_761_dout;
  assign _zz_11057 = _zz_11058;
  assign _zz_11058 = ($signed(_zz_11059) >>> _zz_1523);
  assign _zz_11059 = _zz_11060;
  assign _zz_11060 = ($signed(data_mid_92_real) - $signed(_zz_1521));
  assign _zz_11061 = _zz_11062;
  assign _zz_11062 = ($signed(_zz_11063) >>> _zz_1523);
  assign _zz_11063 = _zz_11064;
  assign _zz_11064 = ($signed(data_mid_92_imag) - $signed(_zz_1522));
  assign _zz_11065 = _zz_11066;
  assign _zz_11066 = ($signed(_zz_11067) >>> _zz_1524);
  assign _zz_11067 = _zz_11068;
  assign _zz_11068 = ($signed(data_mid_92_real) + $signed(_zz_1521));
  assign _zz_11069 = _zz_11070;
  assign _zz_11070 = ($signed(_zz_11071) >>> _zz_1524);
  assign _zz_11071 = _zz_11072;
  assign _zz_11072 = ($signed(data_mid_92_imag) + $signed(_zz_1522));
  assign _zz_11073 = ($signed(twiddle_factor_table_60_real) * $signed(data_mid_125_real));
  assign _zz_11074 = ($signed(twiddle_factor_table_60_imag) * $signed(data_mid_125_imag));
  assign _zz_11075 = fixTo_762_dout;
  assign _zz_11076 = ($signed(twiddle_factor_table_60_real) * $signed(data_mid_125_imag));
  assign _zz_11077 = ($signed(twiddle_factor_table_60_imag) * $signed(data_mid_125_real));
  assign _zz_11078 = fixTo_763_dout;
  assign _zz_11079 = _zz_11080;
  assign _zz_11080 = ($signed(_zz_11081) >>> _zz_1527);
  assign _zz_11081 = _zz_11082;
  assign _zz_11082 = ($signed(data_mid_93_real) - $signed(_zz_1525));
  assign _zz_11083 = _zz_11084;
  assign _zz_11084 = ($signed(_zz_11085) >>> _zz_1527);
  assign _zz_11085 = _zz_11086;
  assign _zz_11086 = ($signed(data_mid_93_imag) - $signed(_zz_1526));
  assign _zz_11087 = _zz_11088;
  assign _zz_11088 = ($signed(_zz_11089) >>> _zz_1528);
  assign _zz_11089 = _zz_11090;
  assign _zz_11090 = ($signed(data_mid_93_real) + $signed(_zz_1525));
  assign _zz_11091 = _zz_11092;
  assign _zz_11092 = ($signed(_zz_11093) >>> _zz_1528);
  assign _zz_11093 = _zz_11094;
  assign _zz_11094 = ($signed(data_mid_93_imag) + $signed(_zz_1526));
  assign _zz_11095 = ($signed(twiddle_factor_table_61_real) * $signed(data_mid_126_real));
  assign _zz_11096 = ($signed(twiddle_factor_table_61_imag) * $signed(data_mid_126_imag));
  assign _zz_11097 = fixTo_764_dout;
  assign _zz_11098 = ($signed(twiddle_factor_table_61_real) * $signed(data_mid_126_imag));
  assign _zz_11099 = ($signed(twiddle_factor_table_61_imag) * $signed(data_mid_126_real));
  assign _zz_11100 = fixTo_765_dout;
  assign _zz_11101 = _zz_11102;
  assign _zz_11102 = ($signed(_zz_11103) >>> _zz_1531);
  assign _zz_11103 = _zz_11104;
  assign _zz_11104 = ($signed(data_mid_94_real) - $signed(_zz_1529));
  assign _zz_11105 = _zz_11106;
  assign _zz_11106 = ($signed(_zz_11107) >>> _zz_1531);
  assign _zz_11107 = _zz_11108;
  assign _zz_11108 = ($signed(data_mid_94_imag) - $signed(_zz_1530));
  assign _zz_11109 = _zz_11110;
  assign _zz_11110 = ($signed(_zz_11111) >>> _zz_1532);
  assign _zz_11111 = _zz_11112;
  assign _zz_11112 = ($signed(data_mid_94_real) + $signed(_zz_1529));
  assign _zz_11113 = _zz_11114;
  assign _zz_11114 = ($signed(_zz_11115) >>> _zz_1532);
  assign _zz_11115 = _zz_11116;
  assign _zz_11116 = ($signed(data_mid_94_imag) + $signed(_zz_1530));
  assign _zz_11117 = ($signed(twiddle_factor_table_62_real) * $signed(data_mid_127_real));
  assign _zz_11118 = ($signed(twiddle_factor_table_62_imag) * $signed(data_mid_127_imag));
  assign _zz_11119 = fixTo_766_dout;
  assign _zz_11120 = ($signed(twiddle_factor_table_62_real) * $signed(data_mid_127_imag));
  assign _zz_11121 = ($signed(twiddle_factor_table_62_imag) * $signed(data_mid_127_real));
  assign _zz_11122 = fixTo_767_dout;
  assign _zz_11123 = _zz_11124;
  assign _zz_11124 = ($signed(_zz_11125) >>> _zz_1535);
  assign _zz_11125 = _zz_11126;
  assign _zz_11126 = ($signed(data_mid_95_real) - $signed(_zz_1533));
  assign _zz_11127 = _zz_11128;
  assign _zz_11128 = ($signed(_zz_11129) >>> _zz_1535);
  assign _zz_11129 = _zz_11130;
  assign _zz_11130 = ($signed(data_mid_95_imag) - $signed(_zz_1534));
  assign _zz_11131 = _zz_11132;
  assign _zz_11132 = ($signed(_zz_11133) >>> _zz_1536);
  assign _zz_11133 = _zz_11134;
  assign _zz_11134 = ($signed(data_mid_95_real) + $signed(_zz_1533));
  assign _zz_11135 = _zz_11136;
  assign _zz_11136 = ($signed(_zz_11137) >>> _zz_1536);
  assign _zz_11137 = _zz_11138;
  assign _zz_11138 = ($signed(data_mid_95_imag) + $signed(_zz_1534));
  assign _zz_11139 = ($signed(twiddle_factor_table_63_real) * $signed(data_mid_64_real));
  assign _zz_11140 = ($signed(twiddle_factor_table_63_imag) * $signed(data_mid_64_imag));
  assign _zz_11141 = fixTo_768_dout;
  assign _zz_11142 = ($signed(twiddle_factor_table_63_real) * $signed(data_mid_64_imag));
  assign _zz_11143 = ($signed(twiddle_factor_table_63_imag) * $signed(data_mid_64_real));
  assign _zz_11144 = fixTo_769_dout;
  assign _zz_11145 = _zz_11146;
  assign _zz_11146 = ($signed(_zz_11147) >>> _zz_1539);
  assign _zz_11147 = _zz_11148;
  assign _zz_11148 = ($signed(data_mid_0_real) - $signed(_zz_1537));
  assign _zz_11149 = _zz_11150;
  assign _zz_11150 = ($signed(_zz_11151) >>> _zz_1539);
  assign _zz_11151 = _zz_11152;
  assign _zz_11152 = ($signed(data_mid_0_imag) - $signed(_zz_1538));
  assign _zz_11153 = _zz_11154;
  assign _zz_11154 = ($signed(_zz_11155) >>> _zz_1540);
  assign _zz_11155 = _zz_11156;
  assign _zz_11156 = ($signed(data_mid_0_real) + $signed(_zz_1537));
  assign _zz_11157 = _zz_11158;
  assign _zz_11158 = ($signed(_zz_11159) >>> _zz_1540);
  assign _zz_11159 = _zz_11160;
  assign _zz_11160 = ($signed(data_mid_0_imag) + $signed(_zz_1538));
  assign _zz_11161 = ($signed(twiddle_factor_table_64_real) * $signed(data_mid_65_real));
  assign _zz_11162 = ($signed(twiddle_factor_table_64_imag) * $signed(data_mid_65_imag));
  assign _zz_11163 = fixTo_770_dout;
  assign _zz_11164 = ($signed(twiddle_factor_table_64_real) * $signed(data_mid_65_imag));
  assign _zz_11165 = ($signed(twiddle_factor_table_64_imag) * $signed(data_mid_65_real));
  assign _zz_11166 = fixTo_771_dout;
  assign _zz_11167 = _zz_11168;
  assign _zz_11168 = ($signed(_zz_11169) >>> _zz_1543);
  assign _zz_11169 = _zz_11170;
  assign _zz_11170 = ($signed(data_mid_1_real) - $signed(_zz_1541));
  assign _zz_11171 = _zz_11172;
  assign _zz_11172 = ($signed(_zz_11173) >>> _zz_1543);
  assign _zz_11173 = _zz_11174;
  assign _zz_11174 = ($signed(data_mid_1_imag) - $signed(_zz_1542));
  assign _zz_11175 = _zz_11176;
  assign _zz_11176 = ($signed(_zz_11177) >>> _zz_1544);
  assign _zz_11177 = _zz_11178;
  assign _zz_11178 = ($signed(data_mid_1_real) + $signed(_zz_1541));
  assign _zz_11179 = _zz_11180;
  assign _zz_11180 = ($signed(_zz_11181) >>> _zz_1544);
  assign _zz_11181 = _zz_11182;
  assign _zz_11182 = ($signed(data_mid_1_imag) + $signed(_zz_1542));
  assign _zz_11183 = ($signed(twiddle_factor_table_65_real) * $signed(data_mid_66_real));
  assign _zz_11184 = ($signed(twiddle_factor_table_65_imag) * $signed(data_mid_66_imag));
  assign _zz_11185 = fixTo_772_dout;
  assign _zz_11186 = ($signed(twiddle_factor_table_65_real) * $signed(data_mid_66_imag));
  assign _zz_11187 = ($signed(twiddle_factor_table_65_imag) * $signed(data_mid_66_real));
  assign _zz_11188 = fixTo_773_dout;
  assign _zz_11189 = _zz_11190;
  assign _zz_11190 = ($signed(_zz_11191) >>> _zz_1547);
  assign _zz_11191 = _zz_11192;
  assign _zz_11192 = ($signed(data_mid_2_real) - $signed(_zz_1545));
  assign _zz_11193 = _zz_11194;
  assign _zz_11194 = ($signed(_zz_11195) >>> _zz_1547);
  assign _zz_11195 = _zz_11196;
  assign _zz_11196 = ($signed(data_mid_2_imag) - $signed(_zz_1546));
  assign _zz_11197 = _zz_11198;
  assign _zz_11198 = ($signed(_zz_11199) >>> _zz_1548);
  assign _zz_11199 = _zz_11200;
  assign _zz_11200 = ($signed(data_mid_2_real) + $signed(_zz_1545));
  assign _zz_11201 = _zz_11202;
  assign _zz_11202 = ($signed(_zz_11203) >>> _zz_1548);
  assign _zz_11203 = _zz_11204;
  assign _zz_11204 = ($signed(data_mid_2_imag) + $signed(_zz_1546));
  assign _zz_11205 = ($signed(twiddle_factor_table_66_real) * $signed(data_mid_67_real));
  assign _zz_11206 = ($signed(twiddle_factor_table_66_imag) * $signed(data_mid_67_imag));
  assign _zz_11207 = fixTo_774_dout;
  assign _zz_11208 = ($signed(twiddle_factor_table_66_real) * $signed(data_mid_67_imag));
  assign _zz_11209 = ($signed(twiddle_factor_table_66_imag) * $signed(data_mid_67_real));
  assign _zz_11210 = fixTo_775_dout;
  assign _zz_11211 = _zz_11212;
  assign _zz_11212 = ($signed(_zz_11213) >>> _zz_1551);
  assign _zz_11213 = _zz_11214;
  assign _zz_11214 = ($signed(data_mid_3_real) - $signed(_zz_1549));
  assign _zz_11215 = _zz_11216;
  assign _zz_11216 = ($signed(_zz_11217) >>> _zz_1551);
  assign _zz_11217 = _zz_11218;
  assign _zz_11218 = ($signed(data_mid_3_imag) - $signed(_zz_1550));
  assign _zz_11219 = _zz_11220;
  assign _zz_11220 = ($signed(_zz_11221) >>> _zz_1552);
  assign _zz_11221 = _zz_11222;
  assign _zz_11222 = ($signed(data_mid_3_real) + $signed(_zz_1549));
  assign _zz_11223 = _zz_11224;
  assign _zz_11224 = ($signed(_zz_11225) >>> _zz_1552);
  assign _zz_11225 = _zz_11226;
  assign _zz_11226 = ($signed(data_mid_3_imag) + $signed(_zz_1550));
  assign _zz_11227 = ($signed(twiddle_factor_table_67_real) * $signed(data_mid_68_real));
  assign _zz_11228 = ($signed(twiddle_factor_table_67_imag) * $signed(data_mid_68_imag));
  assign _zz_11229 = fixTo_776_dout;
  assign _zz_11230 = ($signed(twiddle_factor_table_67_real) * $signed(data_mid_68_imag));
  assign _zz_11231 = ($signed(twiddle_factor_table_67_imag) * $signed(data_mid_68_real));
  assign _zz_11232 = fixTo_777_dout;
  assign _zz_11233 = _zz_11234;
  assign _zz_11234 = ($signed(_zz_11235) >>> _zz_1555);
  assign _zz_11235 = _zz_11236;
  assign _zz_11236 = ($signed(data_mid_4_real) - $signed(_zz_1553));
  assign _zz_11237 = _zz_11238;
  assign _zz_11238 = ($signed(_zz_11239) >>> _zz_1555);
  assign _zz_11239 = _zz_11240;
  assign _zz_11240 = ($signed(data_mid_4_imag) - $signed(_zz_1554));
  assign _zz_11241 = _zz_11242;
  assign _zz_11242 = ($signed(_zz_11243) >>> _zz_1556);
  assign _zz_11243 = _zz_11244;
  assign _zz_11244 = ($signed(data_mid_4_real) + $signed(_zz_1553));
  assign _zz_11245 = _zz_11246;
  assign _zz_11246 = ($signed(_zz_11247) >>> _zz_1556);
  assign _zz_11247 = _zz_11248;
  assign _zz_11248 = ($signed(data_mid_4_imag) + $signed(_zz_1554));
  assign _zz_11249 = ($signed(twiddle_factor_table_68_real) * $signed(data_mid_69_real));
  assign _zz_11250 = ($signed(twiddle_factor_table_68_imag) * $signed(data_mid_69_imag));
  assign _zz_11251 = fixTo_778_dout;
  assign _zz_11252 = ($signed(twiddle_factor_table_68_real) * $signed(data_mid_69_imag));
  assign _zz_11253 = ($signed(twiddle_factor_table_68_imag) * $signed(data_mid_69_real));
  assign _zz_11254 = fixTo_779_dout;
  assign _zz_11255 = _zz_11256;
  assign _zz_11256 = ($signed(_zz_11257) >>> _zz_1559);
  assign _zz_11257 = _zz_11258;
  assign _zz_11258 = ($signed(data_mid_5_real) - $signed(_zz_1557));
  assign _zz_11259 = _zz_11260;
  assign _zz_11260 = ($signed(_zz_11261) >>> _zz_1559);
  assign _zz_11261 = _zz_11262;
  assign _zz_11262 = ($signed(data_mid_5_imag) - $signed(_zz_1558));
  assign _zz_11263 = _zz_11264;
  assign _zz_11264 = ($signed(_zz_11265) >>> _zz_1560);
  assign _zz_11265 = _zz_11266;
  assign _zz_11266 = ($signed(data_mid_5_real) + $signed(_zz_1557));
  assign _zz_11267 = _zz_11268;
  assign _zz_11268 = ($signed(_zz_11269) >>> _zz_1560);
  assign _zz_11269 = _zz_11270;
  assign _zz_11270 = ($signed(data_mid_5_imag) + $signed(_zz_1558));
  assign _zz_11271 = ($signed(twiddle_factor_table_69_real) * $signed(data_mid_70_real));
  assign _zz_11272 = ($signed(twiddle_factor_table_69_imag) * $signed(data_mid_70_imag));
  assign _zz_11273 = fixTo_780_dout;
  assign _zz_11274 = ($signed(twiddle_factor_table_69_real) * $signed(data_mid_70_imag));
  assign _zz_11275 = ($signed(twiddle_factor_table_69_imag) * $signed(data_mid_70_real));
  assign _zz_11276 = fixTo_781_dout;
  assign _zz_11277 = _zz_11278;
  assign _zz_11278 = ($signed(_zz_11279) >>> _zz_1563);
  assign _zz_11279 = _zz_11280;
  assign _zz_11280 = ($signed(data_mid_6_real) - $signed(_zz_1561));
  assign _zz_11281 = _zz_11282;
  assign _zz_11282 = ($signed(_zz_11283) >>> _zz_1563);
  assign _zz_11283 = _zz_11284;
  assign _zz_11284 = ($signed(data_mid_6_imag) - $signed(_zz_1562));
  assign _zz_11285 = _zz_11286;
  assign _zz_11286 = ($signed(_zz_11287) >>> _zz_1564);
  assign _zz_11287 = _zz_11288;
  assign _zz_11288 = ($signed(data_mid_6_real) + $signed(_zz_1561));
  assign _zz_11289 = _zz_11290;
  assign _zz_11290 = ($signed(_zz_11291) >>> _zz_1564);
  assign _zz_11291 = _zz_11292;
  assign _zz_11292 = ($signed(data_mid_6_imag) + $signed(_zz_1562));
  assign _zz_11293 = ($signed(twiddle_factor_table_70_real) * $signed(data_mid_71_real));
  assign _zz_11294 = ($signed(twiddle_factor_table_70_imag) * $signed(data_mid_71_imag));
  assign _zz_11295 = fixTo_782_dout;
  assign _zz_11296 = ($signed(twiddle_factor_table_70_real) * $signed(data_mid_71_imag));
  assign _zz_11297 = ($signed(twiddle_factor_table_70_imag) * $signed(data_mid_71_real));
  assign _zz_11298 = fixTo_783_dout;
  assign _zz_11299 = _zz_11300;
  assign _zz_11300 = ($signed(_zz_11301) >>> _zz_1567);
  assign _zz_11301 = _zz_11302;
  assign _zz_11302 = ($signed(data_mid_7_real) - $signed(_zz_1565));
  assign _zz_11303 = _zz_11304;
  assign _zz_11304 = ($signed(_zz_11305) >>> _zz_1567);
  assign _zz_11305 = _zz_11306;
  assign _zz_11306 = ($signed(data_mid_7_imag) - $signed(_zz_1566));
  assign _zz_11307 = _zz_11308;
  assign _zz_11308 = ($signed(_zz_11309) >>> _zz_1568);
  assign _zz_11309 = _zz_11310;
  assign _zz_11310 = ($signed(data_mid_7_real) + $signed(_zz_1565));
  assign _zz_11311 = _zz_11312;
  assign _zz_11312 = ($signed(_zz_11313) >>> _zz_1568);
  assign _zz_11313 = _zz_11314;
  assign _zz_11314 = ($signed(data_mid_7_imag) + $signed(_zz_1566));
  assign _zz_11315 = ($signed(twiddle_factor_table_71_real) * $signed(data_mid_72_real));
  assign _zz_11316 = ($signed(twiddle_factor_table_71_imag) * $signed(data_mid_72_imag));
  assign _zz_11317 = fixTo_784_dout;
  assign _zz_11318 = ($signed(twiddle_factor_table_71_real) * $signed(data_mid_72_imag));
  assign _zz_11319 = ($signed(twiddle_factor_table_71_imag) * $signed(data_mid_72_real));
  assign _zz_11320 = fixTo_785_dout;
  assign _zz_11321 = _zz_11322;
  assign _zz_11322 = ($signed(_zz_11323) >>> _zz_1571);
  assign _zz_11323 = _zz_11324;
  assign _zz_11324 = ($signed(data_mid_8_real) - $signed(_zz_1569));
  assign _zz_11325 = _zz_11326;
  assign _zz_11326 = ($signed(_zz_11327) >>> _zz_1571);
  assign _zz_11327 = _zz_11328;
  assign _zz_11328 = ($signed(data_mid_8_imag) - $signed(_zz_1570));
  assign _zz_11329 = _zz_11330;
  assign _zz_11330 = ($signed(_zz_11331) >>> _zz_1572);
  assign _zz_11331 = _zz_11332;
  assign _zz_11332 = ($signed(data_mid_8_real) + $signed(_zz_1569));
  assign _zz_11333 = _zz_11334;
  assign _zz_11334 = ($signed(_zz_11335) >>> _zz_1572);
  assign _zz_11335 = _zz_11336;
  assign _zz_11336 = ($signed(data_mid_8_imag) + $signed(_zz_1570));
  assign _zz_11337 = ($signed(twiddle_factor_table_72_real) * $signed(data_mid_73_real));
  assign _zz_11338 = ($signed(twiddle_factor_table_72_imag) * $signed(data_mid_73_imag));
  assign _zz_11339 = fixTo_786_dout;
  assign _zz_11340 = ($signed(twiddle_factor_table_72_real) * $signed(data_mid_73_imag));
  assign _zz_11341 = ($signed(twiddle_factor_table_72_imag) * $signed(data_mid_73_real));
  assign _zz_11342 = fixTo_787_dout;
  assign _zz_11343 = _zz_11344;
  assign _zz_11344 = ($signed(_zz_11345) >>> _zz_1575);
  assign _zz_11345 = _zz_11346;
  assign _zz_11346 = ($signed(data_mid_9_real) - $signed(_zz_1573));
  assign _zz_11347 = _zz_11348;
  assign _zz_11348 = ($signed(_zz_11349) >>> _zz_1575);
  assign _zz_11349 = _zz_11350;
  assign _zz_11350 = ($signed(data_mid_9_imag) - $signed(_zz_1574));
  assign _zz_11351 = _zz_11352;
  assign _zz_11352 = ($signed(_zz_11353) >>> _zz_1576);
  assign _zz_11353 = _zz_11354;
  assign _zz_11354 = ($signed(data_mid_9_real) + $signed(_zz_1573));
  assign _zz_11355 = _zz_11356;
  assign _zz_11356 = ($signed(_zz_11357) >>> _zz_1576);
  assign _zz_11357 = _zz_11358;
  assign _zz_11358 = ($signed(data_mid_9_imag) + $signed(_zz_1574));
  assign _zz_11359 = ($signed(twiddle_factor_table_73_real) * $signed(data_mid_74_real));
  assign _zz_11360 = ($signed(twiddle_factor_table_73_imag) * $signed(data_mid_74_imag));
  assign _zz_11361 = fixTo_788_dout;
  assign _zz_11362 = ($signed(twiddle_factor_table_73_real) * $signed(data_mid_74_imag));
  assign _zz_11363 = ($signed(twiddle_factor_table_73_imag) * $signed(data_mid_74_real));
  assign _zz_11364 = fixTo_789_dout;
  assign _zz_11365 = _zz_11366;
  assign _zz_11366 = ($signed(_zz_11367) >>> _zz_1579);
  assign _zz_11367 = _zz_11368;
  assign _zz_11368 = ($signed(data_mid_10_real) - $signed(_zz_1577));
  assign _zz_11369 = _zz_11370;
  assign _zz_11370 = ($signed(_zz_11371) >>> _zz_1579);
  assign _zz_11371 = _zz_11372;
  assign _zz_11372 = ($signed(data_mid_10_imag) - $signed(_zz_1578));
  assign _zz_11373 = _zz_11374;
  assign _zz_11374 = ($signed(_zz_11375) >>> _zz_1580);
  assign _zz_11375 = _zz_11376;
  assign _zz_11376 = ($signed(data_mid_10_real) + $signed(_zz_1577));
  assign _zz_11377 = _zz_11378;
  assign _zz_11378 = ($signed(_zz_11379) >>> _zz_1580);
  assign _zz_11379 = _zz_11380;
  assign _zz_11380 = ($signed(data_mid_10_imag) + $signed(_zz_1578));
  assign _zz_11381 = ($signed(twiddle_factor_table_74_real) * $signed(data_mid_75_real));
  assign _zz_11382 = ($signed(twiddle_factor_table_74_imag) * $signed(data_mid_75_imag));
  assign _zz_11383 = fixTo_790_dout;
  assign _zz_11384 = ($signed(twiddle_factor_table_74_real) * $signed(data_mid_75_imag));
  assign _zz_11385 = ($signed(twiddle_factor_table_74_imag) * $signed(data_mid_75_real));
  assign _zz_11386 = fixTo_791_dout;
  assign _zz_11387 = _zz_11388;
  assign _zz_11388 = ($signed(_zz_11389) >>> _zz_1583);
  assign _zz_11389 = _zz_11390;
  assign _zz_11390 = ($signed(data_mid_11_real) - $signed(_zz_1581));
  assign _zz_11391 = _zz_11392;
  assign _zz_11392 = ($signed(_zz_11393) >>> _zz_1583);
  assign _zz_11393 = _zz_11394;
  assign _zz_11394 = ($signed(data_mid_11_imag) - $signed(_zz_1582));
  assign _zz_11395 = _zz_11396;
  assign _zz_11396 = ($signed(_zz_11397) >>> _zz_1584);
  assign _zz_11397 = _zz_11398;
  assign _zz_11398 = ($signed(data_mid_11_real) + $signed(_zz_1581));
  assign _zz_11399 = _zz_11400;
  assign _zz_11400 = ($signed(_zz_11401) >>> _zz_1584);
  assign _zz_11401 = _zz_11402;
  assign _zz_11402 = ($signed(data_mid_11_imag) + $signed(_zz_1582));
  assign _zz_11403 = ($signed(twiddle_factor_table_75_real) * $signed(data_mid_76_real));
  assign _zz_11404 = ($signed(twiddle_factor_table_75_imag) * $signed(data_mid_76_imag));
  assign _zz_11405 = fixTo_792_dout;
  assign _zz_11406 = ($signed(twiddle_factor_table_75_real) * $signed(data_mid_76_imag));
  assign _zz_11407 = ($signed(twiddle_factor_table_75_imag) * $signed(data_mid_76_real));
  assign _zz_11408 = fixTo_793_dout;
  assign _zz_11409 = _zz_11410;
  assign _zz_11410 = ($signed(_zz_11411) >>> _zz_1587);
  assign _zz_11411 = _zz_11412;
  assign _zz_11412 = ($signed(data_mid_12_real) - $signed(_zz_1585));
  assign _zz_11413 = _zz_11414;
  assign _zz_11414 = ($signed(_zz_11415) >>> _zz_1587);
  assign _zz_11415 = _zz_11416;
  assign _zz_11416 = ($signed(data_mid_12_imag) - $signed(_zz_1586));
  assign _zz_11417 = _zz_11418;
  assign _zz_11418 = ($signed(_zz_11419) >>> _zz_1588);
  assign _zz_11419 = _zz_11420;
  assign _zz_11420 = ($signed(data_mid_12_real) + $signed(_zz_1585));
  assign _zz_11421 = _zz_11422;
  assign _zz_11422 = ($signed(_zz_11423) >>> _zz_1588);
  assign _zz_11423 = _zz_11424;
  assign _zz_11424 = ($signed(data_mid_12_imag) + $signed(_zz_1586));
  assign _zz_11425 = ($signed(twiddle_factor_table_76_real) * $signed(data_mid_77_real));
  assign _zz_11426 = ($signed(twiddle_factor_table_76_imag) * $signed(data_mid_77_imag));
  assign _zz_11427 = fixTo_794_dout;
  assign _zz_11428 = ($signed(twiddle_factor_table_76_real) * $signed(data_mid_77_imag));
  assign _zz_11429 = ($signed(twiddle_factor_table_76_imag) * $signed(data_mid_77_real));
  assign _zz_11430 = fixTo_795_dout;
  assign _zz_11431 = _zz_11432;
  assign _zz_11432 = ($signed(_zz_11433) >>> _zz_1591);
  assign _zz_11433 = _zz_11434;
  assign _zz_11434 = ($signed(data_mid_13_real) - $signed(_zz_1589));
  assign _zz_11435 = _zz_11436;
  assign _zz_11436 = ($signed(_zz_11437) >>> _zz_1591);
  assign _zz_11437 = _zz_11438;
  assign _zz_11438 = ($signed(data_mid_13_imag) - $signed(_zz_1590));
  assign _zz_11439 = _zz_11440;
  assign _zz_11440 = ($signed(_zz_11441) >>> _zz_1592);
  assign _zz_11441 = _zz_11442;
  assign _zz_11442 = ($signed(data_mid_13_real) + $signed(_zz_1589));
  assign _zz_11443 = _zz_11444;
  assign _zz_11444 = ($signed(_zz_11445) >>> _zz_1592);
  assign _zz_11445 = _zz_11446;
  assign _zz_11446 = ($signed(data_mid_13_imag) + $signed(_zz_1590));
  assign _zz_11447 = ($signed(twiddle_factor_table_77_real) * $signed(data_mid_78_real));
  assign _zz_11448 = ($signed(twiddle_factor_table_77_imag) * $signed(data_mid_78_imag));
  assign _zz_11449 = fixTo_796_dout;
  assign _zz_11450 = ($signed(twiddle_factor_table_77_real) * $signed(data_mid_78_imag));
  assign _zz_11451 = ($signed(twiddle_factor_table_77_imag) * $signed(data_mid_78_real));
  assign _zz_11452 = fixTo_797_dout;
  assign _zz_11453 = _zz_11454;
  assign _zz_11454 = ($signed(_zz_11455) >>> _zz_1595);
  assign _zz_11455 = _zz_11456;
  assign _zz_11456 = ($signed(data_mid_14_real) - $signed(_zz_1593));
  assign _zz_11457 = _zz_11458;
  assign _zz_11458 = ($signed(_zz_11459) >>> _zz_1595);
  assign _zz_11459 = _zz_11460;
  assign _zz_11460 = ($signed(data_mid_14_imag) - $signed(_zz_1594));
  assign _zz_11461 = _zz_11462;
  assign _zz_11462 = ($signed(_zz_11463) >>> _zz_1596);
  assign _zz_11463 = _zz_11464;
  assign _zz_11464 = ($signed(data_mid_14_real) + $signed(_zz_1593));
  assign _zz_11465 = _zz_11466;
  assign _zz_11466 = ($signed(_zz_11467) >>> _zz_1596);
  assign _zz_11467 = _zz_11468;
  assign _zz_11468 = ($signed(data_mid_14_imag) + $signed(_zz_1594));
  assign _zz_11469 = ($signed(twiddle_factor_table_78_real) * $signed(data_mid_79_real));
  assign _zz_11470 = ($signed(twiddle_factor_table_78_imag) * $signed(data_mid_79_imag));
  assign _zz_11471 = fixTo_798_dout;
  assign _zz_11472 = ($signed(twiddle_factor_table_78_real) * $signed(data_mid_79_imag));
  assign _zz_11473 = ($signed(twiddle_factor_table_78_imag) * $signed(data_mid_79_real));
  assign _zz_11474 = fixTo_799_dout;
  assign _zz_11475 = _zz_11476;
  assign _zz_11476 = ($signed(_zz_11477) >>> _zz_1599);
  assign _zz_11477 = _zz_11478;
  assign _zz_11478 = ($signed(data_mid_15_real) - $signed(_zz_1597));
  assign _zz_11479 = _zz_11480;
  assign _zz_11480 = ($signed(_zz_11481) >>> _zz_1599);
  assign _zz_11481 = _zz_11482;
  assign _zz_11482 = ($signed(data_mid_15_imag) - $signed(_zz_1598));
  assign _zz_11483 = _zz_11484;
  assign _zz_11484 = ($signed(_zz_11485) >>> _zz_1600);
  assign _zz_11485 = _zz_11486;
  assign _zz_11486 = ($signed(data_mid_15_real) + $signed(_zz_1597));
  assign _zz_11487 = _zz_11488;
  assign _zz_11488 = ($signed(_zz_11489) >>> _zz_1600);
  assign _zz_11489 = _zz_11490;
  assign _zz_11490 = ($signed(data_mid_15_imag) + $signed(_zz_1598));
  assign _zz_11491 = ($signed(twiddle_factor_table_79_real) * $signed(data_mid_80_real));
  assign _zz_11492 = ($signed(twiddle_factor_table_79_imag) * $signed(data_mid_80_imag));
  assign _zz_11493 = fixTo_800_dout;
  assign _zz_11494 = ($signed(twiddle_factor_table_79_real) * $signed(data_mid_80_imag));
  assign _zz_11495 = ($signed(twiddle_factor_table_79_imag) * $signed(data_mid_80_real));
  assign _zz_11496 = fixTo_801_dout;
  assign _zz_11497 = _zz_11498;
  assign _zz_11498 = ($signed(_zz_11499) >>> _zz_1603);
  assign _zz_11499 = _zz_11500;
  assign _zz_11500 = ($signed(data_mid_16_real) - $signed(_zz_1601));
  assign _zz_11501 = _zz_11502;
  assign _zz_11502 = ($signed(_zz_11503) >>> _zz_1603);
  assign _zz_11503 = _zz_11504;
  assign _zz_11504 = ($signed(data_mid_16_imag) - $signed(_zz_1602));
  assign _zz_11505 = _zz_11506;
  assign _zz_11506 = ($signed(_zz_11507) >>> _zz_1604);
  assign _zz_11507 = _zz_11508;
  assign _zz_11508 = ($signed(data_mid_16_real) + $signed(_zz_1601));
  assign _zz_11509 = _zz_11510;
  assign _zz_11510 = ($signed(_zz_11511) >>> _zz_1604);
  assign _zz_11511 = _zz_11512;
  assign _zz_11512 = ($signed(data_mid_16_imag) + $signed(_zz_1602));
  assign _zz_11513 = ($signed(twiddle_factor_table_80_real) * $signed(data_mid_81_real));
  assign _zz_11514 = ($signed(twiddle_factor_table_80_imag) * $signed(data_mid_81_imag));
  assign _zz_11515 = fixTo_802_dout;
  assign _zz_11516 = ($signed(twiddle_factor_table_80_real) * $signed(data_mid_81_imag));
  assign _zz_11517 = ($signed(twiddle_factor_table_80_imag) * $signed(data_mid_81_real));
  assign _zz_11518 = fixTo_803_dout;
  assign _zz_11519 = _zz_11520;
  assign _zz_11520 = ($signed(_zz_11521) >>> _zz_1607);
  assign _zz_11521 = _zz_11522;
  assign _zz_11522 = ($signed(data_mid_17_real) - $signed(_zz_1605));
  assign _zz_11523 = _zz_11524;
  assign _zz_11524 = ($signed(_zz_11525) >>> _zz_1607);
  assign _zz_11525 = _zz_11526;
  assign _zz_11526 = ($signed(data_mid_17_imag) - $signed(_zz_1606));
  assign _zz_11527 = _zz_11528;
  assign _zz_11528 = ($signed(_zz_11529) >>> _zz_1608);
  assign _zz_11529 = _zz_11530;
  assign _zz_11530 = ($signed(data_mid_17_real) + $signed(_zz_1605));
  assign _zz_11531 = _zz_11532;
  assign _zz_11532 = ($signed(_zz_11533) >>> _zz_1608);
  assign _zz_11533 = _zz_11534;
  assign _zz_11534 = ($signed(data_mid_17_imag) + $signed(_zz_1606));
  assign _zz_11535 = ($signed(twiddle_factor_table_81_real) * $signed(data_mid_82_real));
  assign _zz_11536 = ($signed(twiddle_factor_table_81_imag) * $signed(data_mid_82_imag));
  assign _zz_11537 = fixTo_804_dout;
  assign _zz_11538 = ($signed(twiddle_factor_table_81_real) * $signed(data_mid_82_imag));
  assign _zz_11539 = ($signed(twiddle_factor_table_81_imag) * $signed(data_mid_82_real));
  assign _zz_11540 = fixTo_805_dout;
  assign _zz_11541 = _zz_11542;
  assign _zz_11542 = ($signed(_zz_11543) >>> _zz_1611);
  assign _zz_11543 = _zz_11544;
  assign _zz_11544 = ($signed(data_mid_18_real) - $signed(_zz_1609));
  assign _zz_11545 = _zz_11546;
  assign _zz_11546 = ($signed(_zz_11547) >>> _zz_1611);
  assign _zz_11547 = _zz_11548;
  assign _zz_11548 = ($signed(data_mid_18_imag) - $signed(_zz_1610));
  assign _zz_11549 = _zz_11550;
  assign _zz_11550 = ($signed(_zz_11551) >>> _zz_1612);
  assign _zz_11551 = _zz_11552;
  assign _zz_11552 = ($signed(data_mid_18_real) + $signed(_zz_1609));
  assign _zz_11553 = _zz_11554;
  assign _zz_11554 = ($signed(_zz_11555) >>> _zz_1612);
  assign _zz_11555 = _zz_11556;
  assign _zz_11556 = ($signed(data_mid_18_imag) + $signed(_zz_1610));
  assign _zz_11557 = ($signed(twiddle_factor_table_82_real) * $signed(data_mid_83_real));
  assign _zz_11558 = ($signed(twiddle_factor_table_82_imag) * $signed(data_mid_83_imag));
  assign _zz_11559 = fixTo_806_dout;
  assign _zz_11560 = ($signed(twiddle_factor_table_82_real) * $signed(data_mid_83_imag));
  assign _zz_11561 = ($signed(twiddle_factor_table_82_imag) * $signed(data_mid_83_real));
  assign _zz_11562 = fixTo_807_dout;
  assign _zz_11563 = _zz_11564;
  assign _zz_11564 = ($signed(_zz_11565) >>> _zz_1615);
  assign _zz_11565 = _zz_11566;
  assign _zz_11566 = ($signed(data_mid_19_real) - $signed(_zz_1613));
  assign _zz_11567 = _zz_11568;
  assign _zz_11568 = ($signed(_zz_11569) >>> _zz_1615);
  assign _zz_11569 = _zz_11570;
  assign _zz_11570 = ($signed(data_mid_19_imag) - $signed(_zz_1614));
  assign _zz_11571 = _zz_11572;
  assign _zz_11572 = ($signed(_zz_11573) >>> _zz_1616);
  assign _zz_11573 = _zz_11574;
  assign _zz_11574 = ($signed(data_mid_19_real) + $signed(_zz_1613));
  assign _zz_11575 = _zz_11576;
  assign _zz_11576 = ($signed(_zz_11577) >>> _zz_1616);
  assign _zz_11577 = _zz_11578;
  assign _zz_11578 = ($signed(data_mid_19_imag) + $signed(_zz_1614));
  assign _zz_11579 = ($signed(twiddle_factor_table_83_real) * $signed(data_mid_84_real));
  assign _zz_11580 = ($signed(twiddle_factor_table_83_imag) * $signed(data_mid_84_imag));
  assign _zz_11581 = fixTo_808_dout;
  assign _zz_11582 = ($signed(twiddle_factor_table_83_real) * $signed(data_mid_84_imag));
  assign _zz_11583 = ($signed(twiddle_factor_table_83_imag) * $signed(data_mid_84_real));
  assign _zz_11584 = fixTo_809_dout;
  assign _zz_11585 = _zz_11586;
  assign _zz_11586 = ($signed(_zz_11587) >>> _zz_1619);
  assign _zz_11587 = _zz_11588;
  assign _zz_11588 = ($signed(data_mid_20_real) - $signed(_zz_1617));
  assign _zz_11589 = _zz_11590;
  assign _zz_11590 = ($signed(_zz_11591) >>> _zz_1619);
  assign _zz_11591 = _zz_11592;
  assign _zz_11592 = ($signed(data_mid_20_imag) - $signed(_zz_1618));
  assign _zz_11593 = _zz_11594;
  assign _zz_11594 = ($signed(_zz_11595) >>> _zz_1620);
  assign _zz_11595 = _zz_11596;
  assign _zz_11596 = ($signed(data_mid_20_real) + $signed(_zz_1617));
  assign _zz_11597 = _zz_11598;
  assign _zz_11598 = ($signed(_zz_11599) >>> _zz_1620);
  assign _zz_11599 = _zz_11600;
  assign _zz_11600 = ($signed(data_mid_20_imag) + $signed(_zz_1618));
  assign _zz_11601 = ($signed(twiddle_factor_table_84_real) * $signed(data_mid_85_real));
  assign _zz_11602 = ($signed(twiddle_factor_table_84_imag) * $signed(data_mid_85_imag));
  assign _zz_11603 = fixTo_810_dout;
  assign _zz_11604 = ($signed(twiddle_factor_table_84_real) * $signed(data_mid_85_imag));
  assign _zz_11605 = ($signed(twiddle_factor_table_84_imag) * $signed(data_mid_85_real));
  assign _zz_11606 = fixTo_811_dout;
  assign _zz_11607 = _zz_11608;
  assign _zz_11608 = ($signed(_zz_11609) >>> _zz_1623);
  assign _zz_11609 = _zz_11610;
  assign _zz_11610 = ($signed(data_mid_21_real) - $signed(_zz_1621));
  assign _zz_11611 = _zz_11612;
  assign _zz_11612 = ($signed(_zz_11613) >>> _zz_1623);
  assign _zz_11613 = _zz_11614;
  assign _zz_11614 = ($signed(data_mid_21_imag) - $signed(_zz_1622));
  assign _zz_11615 = _zz_11616;
  assign _zz_11616 = ($signed(_zz_11617) >>> _zz_1624);
  assign _zz_11617 = _zz_11618;
  assign _zz_11618 = ($signed(data_mid_21_real) + $signed(_zz_1621));
  assign _zz_11619 = _zz_11620;
  assign _zz_11620 = ($signed(_zz_11621) >>> _zz_1624);
  assign _zz_11621 = _zz_11622;
  assign _zz_11622 = ($signed(data_mid_21_imag) + $signed(_zz_1622));
  assign _zz_11623 = ($signed(twiddle_factor_table_85_real) * $signed(data_mid_86_real));
  assign _zz_11624 = ($signed(twiddle_factor_table_85_imag) * $signed(data_mid_86_imag));
  assign _zz_11625 = fixTo_812_dout;
  assign _zz_11626 = ($signed(twiddle_factor_table_85_real) * $signed(data_mid_86_imag));
  assign _zz_11627 = ($signed(twiddle_factor_table_85_imag) * $signed(data_mid_86_real));
  assign _zz_11628 = fixTo_813_dout;
  assign _zz_11629 = _zz_11630;
  assign _zz_11630 = ($signed(_zz_11631) >>> _zz_1627);
  assign _zz_11631 = _zz_11632;
  assign _zz_11632 = ($signed(data_mid_22_real) - $signed(_zz_1625));
  assign _zz_11633 = _zz_11634;
  assign _zz_11634 = ($signed(_zz_11635) >>> _zz_1627);
  assign _zz_11635 = _zz_11636;
  assign _zz_11636 = ($signed(data_mid_22_imag) - $signed(_zz_1626));
  assign _zz_11637 = _zz_11638;
  assign _zz_11638 = ($signed(_zz_11639) >>> _zz_1628);
  assign _zz_11639 = _zz_11640;
  assign _zz_11640 = ($signed(data_mid_22_real) + $signed(_zz_1625));
  assign _zz_11641 = _zz_11642;
  assign _zz_11642 = ($signed(_zz_11643) >>> _zz_1628);
  assign _zz_11643 = _zz_11644;
  assign _zz_11644 = ($signed(data_mid_22_imag) + $signed(_zz_1626));
  assign _zz_11645 = ($signed(twiddle_factor_table_86_real) * $signed(data_mid_87_real));
  assign _zz_11646 = ($signed(twiddle_factor_table_86_imag) * $signed(data_mid_87_imag));
  assign _zz_11647 = fixTo_814_dout;
  assign _zz_11648 = ($signed(twiddle_factor_table_86_real) * $signed(data_mid_87_imag));
  assign _zz_11649 = ($signed(twiddle_factor_table_86_imag) * $signed(data_mid_87_real));
  assign _zz_11650 = fixTo_815_dout;
  assign _zz_11651 = _zz_11652;
  assign _zz_11652 = ($signed(_zz_11653) >>> _zz_1631);
  assign _zz_11653 = _zz_11654;
  assign _zz_11654 = ($signed(data_mid_23_real) - $signed(_zz_1629));
  assign _zz_11655 = _zz_11656;
  assign _zz_11656 = ($signed(_zz_11657) >>> _zz_1631);
  assign _zz_11657 = _zz_11658;
  assign _zz_11658 = ($signed(data_mid_23_imag) - $signed(_zz_1630));
  assign _zz_11659 = _zz_11660;
  assign _zz_11660 = ($signed(_zz_11661) >>> _zz_1632);
  assign _zz_11661 = _zz_11662;
  assign _zz_11662 = ($signed(data_mid_23_real) + $signed(_zz_1629));
  assign _zz_11663 = _zz_11664;
  assign _zz_11664 = ($signed(_zz_11665) >>> _zz_1632);
  assign _zz_11665 = _zz_11666;
  assign _zz_11666 = ($signed(data_mid_23_imag) + $signed(_zz_1630));
  assign _zz_11667 = ($signed(twiddle_factor_table_87_real) * $signed(data_mid_88_real));
  assign _zz_11668 = ($signed(twiddle_factor_table_87_imag) * $signed(data_mid_88_imag));
  assign _zz_11669 = fixTo_816_dout;
  assign _zz_11670 = ($signed(twiddle_factor_table_87_real) * $signed(data_mid_88_imag));
  assign _zz_11671 = ($signed(twiddle_factor_table_87_imag) * $signed(data_mid_88_real));
  assign _zz_11672 = fixTo_817_dout;
  assign _zz_11673 = _zz_11674;
  assign _zz_11674 = ($signed(_zz_11675) >>> _zz_1635);
  assign _zz_11675 = _zz_11676;
  assign _zz_11676 = ($signed(data_mid_24_real) - $signed(_zz_1633));
  assign _zz_11677 = _zz_11678;
  assign _zz_11678 = ($signed(_zz_11679) >>> _zz_1635);
  assign _zz_11679 = _zz_11680;
  assign _zz_11680 = ($signed(data_mid_24_imag) - $signed(_zz_1634));
  assign _zz_11681 = _zz_11682;
  assign _zz_11682 = ($signed(_zz_11683) >>> _zz_1636);
  assign _zz_11683 = _zz_11684;
  assign _zz_11684 = ($signed(data_mid_24_real) + $signed(_zz_1633));
  assign _zz_11685 = _zz_11686;
  assign _zz_11686 = ($signed(_zz_11687) >>> _zz_1636);
  assign _zz_11687 = _zz_11688;
  assign _zz_11688 = ($signed(data_mid_24_imag) + $signed(_zz_1634));
  assign _zz_11689 = ($signed(twiddle_factor_table_88_real) * $signed(data_mid_89_real));
  assign _zz_11690 = ($signed(twiddle_factor_table_88_imag) * $signed(data_mid_89_imag));
  assign _zz_11691 = fixTo_818_dout;
  assign _zz_11692 = ($signed(twiddle_factor_table_88_real) * $signed(data_mid_89_imag));
  assign _zz_11693 = ($signed(twiddle_factor_table_88_imag) * $signed(data_mid_89_real));
  assign _zz_11694 = fixTo_819_dout;
  assign _zz_11695 = _zz_11696;
  assign _zz_11696 = ($signed(_zz_11697) >>> _zz_1639);
  assign _zz_11697 = _zz_11698;
  assign _zz_11698 = ($signed(data_mid_25_real) - $signed(_zz_1637));
  assign _zz_11699 = _zz_11700;
  assign _zz_11700 = ($signed(_zz_11701) >>> _zz_1639);
  assign _zz_11701 = _zz_11702;
  assign _zz_11702 = ($signed(data_mid_25_imag) - $signed(_zz_1638));
  assign _zz_11703 = _zz_11704;
  assign _zz_11704 = ($signed(_zz_11705) >>> _zz_1640);
  assign _zz_11705 = _zz_11706;
  assign _zz_11706 = ($signed(data_mid_25_real) + $signed(_zz_1637));
  assign _zz_11707 = _zz_11708;
  assign _zz_11708 = ($signed(_zz_11709) >>> _zz_1640);
  assign _zz_11709 = _zz_11710;
  assign _zz_11710 = ($signed(data_mid_25_imag) + $signed(_zz_1638));
  assign _zz_11711 = ($signed(twiddle_factor_table_89_real) * $signed(data_mid_90_real));
  assign _zz_11712 = ($signed(twiddle_factor_table_89_imag) * $signed(data_mid_90_imag));
  assign _zz_11713 = fixTo_820_dout;
  assign _zz_11714 = ($signed(twiddle_factor_table_89_real) * $signed(data_mid_90_imag));
  assign _zz_11715 = ($signed(twiddle_factor_table_89_imag) * $signed(data_mid_90_real));
  assign _zz_11716 = fixTo_821_dout;
  assign _zz_11717 = _zz_11718;
  assign _zz_11718 = ($signed(_zz_11719) >>> _zz_1643);
  assign _zz_11719 = _zz_11720;
  assign _zz_11720 = ($signed(data_mid_26_real) - $signed(_zz_1641));
  assign _zz_11721 = _zz_11722;
  assign _zz_11722 = ($signed(_zz_11723) >>> _zz_1643);
  assign _zz_11723 = _zz_11724;
  assign _zz_11724 = ($signed(data_mid_26_imag) - $signed(_zz_1642));
  assign _zz_11725 = _zz_11726;
  assign _zz_11726 = ($signed(_zz_11727) >>> _zz_1644);
  assign _zz_11727 = _zz_11728;
  assign _zz_11728 = ($signed(data_mid_26_real) + $signed(_zz_1641));
  assign _zz_11729 = _zz_11730;
  assign _zz_11730 = ($signed(_zz_11731) >>> _zz_1644);
  assign _zz_11731 = _zz_11732;
  assign _zz_11732 = ($signed(data_mid_26_imag) + $signed(_zz_1642));
  assign _zz_11733 = ($signed(twiddle_factor_table_90_real) * $signed(data_mid_91_real));
  assign _zz_11734 = ($signed(twiddle_factor_table_90_imag) * $signed(data_mid_91_imag));
  assign _zz_11735 = fixTo_822_dout;
  assign _zz_11736 = ($signed(twiddle_factor_table_90_real) * $signed(data_mid_91_imag));
  assign _zz_11737 = ($signed(twiddle_factor_table_90_imag) * $signed(data_mid_91_real));
  assign _zz_11738 = fixTo_823_dout;
  assign _zz_11739 = _zz_11740;
  assign _zz_11740 = ($signed(_zz_11741) >>> _zz_1647);
  assign _zz_11741 = _zz_11742;
  assign _zz_11742 = ($signed(data_mid_27_real) - $signed(_zz_1645));
  assign _zz_11743 = _zz_11744;
  assign _zz_11744 = ($signed(_zz_11745) >>> _zz_1647);
  assign _zz_11745 = _zz_11746;
  assign _zz_11746 = ($signed(data_mid_27_imag) - $signed(_zz_1646));
  assign _zz_11747 = _zz_11748;
  assign _zz_11748 = ($signed(_zz_11749) >>> _zz_1648);
  assign _zz_11749 = _zz_11750;
  assign _zz_11750 = ($signed(data_mid_27_real) + $signed(_zz_1645));
  assign _zz_11751 = _zz_11752;
  assign _zz_11752 = ($signed(_zz_11753) >>> _zz_1648);
  assign _zz_11753 = _zz_11754;
  assign _zz_11754 = ($signed(data_mid_27_imag) + $signed(_zz_1646));
  assign _zz_11755 = ($signed(twiddle_factor_table_91_real) * $signed(data_mid_92_real));
  assign _zz_11756 = ($signed(twiddle_factor_table_91_imag) * $signed(data_mid_92_imag));
  assign _zz_11757 = fixTo_824_dout;
  assign _zz_11758 = ($signed(twiddle_factor_table_91_real) * $signed(data_mid_92_imag));
  assign _zz_11759 = ($signed(twiddle_factor_table_91_imag) * $signed(data_mid_92_real));
  assign _zz_11760 = fixTo_825_dout;
  assign _zz_11761 = _zz_11762;
  assign _zz_11762 = ($signed(_zz_11763) >>> _zz_1651);
  assign _zz_11763 = _zz_11764;
  assign _zz_11764 = ($signed(data_mid_28_real) - $signed(_zz_1649));
  assign _zz_11765 = _zz_11766;
  assign _zz_11766 = ($signed(_zz_11767) >>> _zz_1651);
  assign _zz_11767 = _zz_11768;
  assign _zz_11768 = ($signed(data_mid_28_imag) - $signed(_zz_1650));
  assign _zz_11769 = _zz_11770;
  assign _zz_11770 = ($signed(_zz_11771) >>> _zz_1652);
  assign _zz_11771 = _zz_11772;
  assign _zz_11772 = ($signed(data_mid_28_real) + $signed(_zz_1649));
  assign _zz_11773 = _zz_11774;
  assign _zz_11774 = ($signed(_zz_11775) >>> _zz_1652);
  assign _zz_11775 = _zz_11776;
  assign _zz_11776 = ($signed(data_mid_28_imag) + $signed(_zz_1650));
  assign _zz_11777 = ($signed(twiddle_factor_table_92_real) * $signed(data_mid_93_real));
  assign _zz_11778 = ($signed(twiddle_factor_table_92_imag) * $signed(data_mid_93_imag));
  assign _zz_11779 = fixTo_826_dout;
  assign _zz_11780 = ($signed(twiddle_factor_table_92_real) * $signed(data_mid_93_imag));
  assign _zz_11781 = ($signed(twiddle_factor_table_92_imag) * $signed(data_mid_93_real));
  assign _zz_11782 = fixTo_827_dout;
  assign _zz_11783 = _zz_11784;
  assign _zz_11784 = ($signed(_zz_11785) >>> _zz_1655);
  assign _zz_11785 = _zz_11786;
  assign _zz_11786 = ($signed(data_mid_29_real) - $signed(_zz_1653));
  assign _zz_11787 = _zz_11788;
  assign _zz_11788 = ($signed(_zz_11789) >>> _zz_1655);
  assign _zz_11789 = _zz_11790;
  assign _zz_11790 = ($signed(data_mid_29_imag) - $signed(_zz_1654));
  assign _zz_11791 = _zz_11792;
  assign _zz_11792 = ($signed(_zz_11793) >>> _zz_1656);
  assign _zz_11793 = _zz_11794;
  assign _zz_11794 = ($signed(data_mid_29_real) + $signed(_zz_1653));
  assign _zz_11795 = _zz_11796;
  assign _zz_11796 = ($signed(_zz_11797) >>> _zz_1656);
  assign _zz_11797 = _zz_11798;
  assign _zz_11798 = ($signed(data_mid_29_imag) + $signed(_zz_1654));
  assign _zz_11799 = ($signed(twiddle_factor_table_93_real) * $signed(data_mid_94_real));
  assign _zz_11800 = ($signed(twiddle_factor_table_93_imag) * $signed(data_mid_94_imag));
  assign _zz_11801 = fixTo_828_dout;
  assign _zz_11802 = ($signed(twiddle_factor_table_93_real) * $signed(data_mid_94_imag));
  assign _zz_11803 = ($signed(twiddle_factor_table_93_imag) * $signed(data_mid_94_real));
  assign _zz_11804 = fixTo_829_dout;
  assign _zz_11805 = _zz_11806;
  assign _zz_11806 = ($signed(_zz_11807) >>> _zz_1659);
  assign _zz_11807 = _zz_11808;
  assign _zz_11808 = ($signed(data_mid_30_real) - $signed(_zz_1657));
  assign _zz_11809 = _zz_11810;
  assign _zz_11810 = ($signed(_zz_11811) >>> _zz_1659);
  assign _zz_11811 = _zz_11812;
  assign _zz_11812 = ($signed(data_mid_30_imag) - $signed(_zz_1658));
  assign _zz_11813 = _zz_11814;
  assign _zz_11814 = ($signed(_zz_11815) >>> _zz_1660);
  assign _zz_11815 = _zz_11816;
  assign _zz_11816 = ($signed(data_mid_30_real) + $signed(_zz_1657));
  assign _zz_11817 = _zz_11818;
  assign _zz_11818 = ($signed(_zz_11819) >>> _zz_1660);
  assign _zz_11819 = _zz_11820;
  assign _zz_11820 = ($signed(data_mid_30_imag) + $signed(_zz_1658));
  assign _zz_11821 = ($signed(twiddle_factor_table_94_real) * $signed(data_mid_95_real));
  assign _zz_11822 = ($signed(twiddle_factor_table_94_imag) * $signed(data_mid_95_imag));
  assign _zz_11823 = fixTo_830_dout;
  assign _zz_11824 = ($signed(twiddle_factor_table_94_real) * $signed(data_mid_95_imag));
  assign _zz_11825 = ($signed(twiddle_factor_table_94_imag) * $signed(data_mid_95_real));
  assign _zz_11826 = fixTo_831_dout;
  assign _zz_11827 = _zz_11828;
  assign _zz_11828 = ($signed(_zz_11829) >>> _zz_1663);
  assign _zz_11829 = _zz_11830;
  assign _zz_11830 = ($signed(data_mid_31_real) - $signed(_zz_1661));
  assign _zz_11831 = _zz_11832;
  assign _zz_11832 = ($signed(_zz_11833) >>> _zz_1663);
  assign _zz_11833 = _zz_11834;
  assign _zz_11834 = ($signed(data_mid_31_imag) - $signed(_zz_1662));
  assign _zz_11835 = _zz_11836;
  assign _zz_11836 = ($signed(_zz_11837) >>> _zz_1664);
  assign _zz_11837 = _zz_11838;
  assign _zz_11838 = ($signed(data_mid_31_real) + $signed(_zz_1661));
  assign _zz_11839 = _zz_11840;
  assign _zz_11840 = ($signed(_zz_11841) >>> _zz_1664);
  assign _zz_11841 = _zz_11842;
  assign _zz_11842 = ($signed(data_mid_31_imag) + $signed(_zz_1662));
  assign _zz_11843 = ($signed(twiddle_factor_table_95_real) * $signed(data_mid_96_real));
  assign _zz_11844 = ($signed(twiddle_factor_table_95_imag) * $signed(data_mid_96_imag));
  assign _zz_11845 = fixTo_832_dout;
  assign _zz_11846 = ($signed(twiddle_factor_table_95_real) * $signed(data_mid_96_imag));
  assign _zz_11847 = ($signed(twiddle_factor_table_95_imag) * $signed(data_mid_96_real));
  assign _zz_11848 = fixTo_833_dout;
  assign _zz_11849 = _zz_11850;
  assign _zz_11850 = ($signed(_zz_11851) >>> _zz_1667);
  assign _zz_11851 = _zz_11852;
  assign _zz_11852 = ($signed(data_mid_32_real) - $signed(_zz_1665));
  assign _zz_11853 = _zz_11854;
  assign _zz_11854 = ($signed(_zz_11855) >>> _zz_1667);
  assign _zz_11855 = _zz_11856;
  assign _zz_11856 = ($signed(data_mid_32_imag) - $signed(_zz_1666));
  assign _zz_11857 = _zz_11858;
  assign _zz_11858 = ($signed(_zz_11859) >>> _zz_1668);
  assign _zz_11859 = _zz_11860;
  assign _zz_11860 = ($signed(data_mid_32_real) + $signed(_zz_1665));
  assign _zz_11861 = _zz_11862;
  assign _zz_11862 = ($signed(_zz_11863) >>> _zz_1668);
  assign _zz_11863 = _zz_11864;
  assign _zz_11864 = ($signed(data_mid_32_imag) + $signed(_zz_1666));
  assign _zz_11865 = ($signed(twiddle_factor_table_96_real) * $signed(data_mid_97_real));
  assign _zz_11866 = ($signed(twiddle_factor_table_96_imag) * $signed(data_mid_97_imag));
  assign _zz_11867 = fixTo_834_dout;
  assign _zz_11868 = ($signed(twiddle_factor_table_96_real) * $signed(data_mid_97_imag));
  assign _zz_11869 = ($signed(twiddle_factor_table_96_imag) * $signed(data_mid_97_real));
  assign _zz_11870 = fixTo_835_dout;
  assign _zz_11871 = _zz_11872;
  assign _zz_11872 = ($signed(_zz_11873) >>> _zz_1671);
  assign _zz_11873 = _zz_11874;
  assign _zz_11874 = ($signed(data_mid_33_real) - $signed(_zz_1669));
  assign _zz_11875 = _zz_11876;
  assign _zz_11876 = ($signed(_zz_11877) >>> _zz_1671);
  assign _zz_11877 = _zz_11878;
  assign _zz_11878 = ($signed(data_mid_33_imag) - $signed(_zz_1670));
  assign _zz_11879 = _zz_11880;
  assign _zz_11880 = ($signed(_zz_11881) >>> _zz_1672);
  assign _zz_11881 = _zz_11882;
  assign _zz_11882 = ($signed(data_mid_33_real) + $signed(_zz_1669));
  assign _zz_11883 = _zz_11884;
  assign _zz_11884 = ($signed(_zz_11885) >>> _zz_1672);
  assign _zz_11885 = _zz_11886;
  assign _zz_11886 = ($signed(data_mid_33_imag) + $signed(_zz_1670));
  assign _zz_11887 = ($signed(twiddle_factor_table_97_real) * $signed(data_mid_98_real));
  assign _zz_11888 = ($signed(twiddle_factor_table_97_imag) * $signed(data_mid_98_imag));
  assign _zz_11889 = fixTo_836_dout;
  assign _zz_11890 = ($signed(twiddle_factor_table_97_real) * $signed(data_mid_98_imag));
  assign _zz_11891 = ($signed(twiddle_factor_table_97_imag) * $signed(data_mid_98_real));
  assign _zz_11892 = fixTo_837_dout;
  assign _zz_11893 = _zz_11894;
  assign _zz_11894 = ($signed(_zz_11895) >>> _zz_1675);
  assign _zz_11895 = _zz_11896;
  assign _zz_11896 = ($signed(data_mid_34_real) - $signed(_zz_1673));
  assign _zz_11897 = _zz_11898;
  assign _zz_11898 = ($signed(_zz_11899) >>> _zz_1675);
  assign _zz_11899 = _zz_11900;
  assign _zz_11900 = ($signed(data_mid_34_imag) - $signed(_zz_1674));
  assign _zz_11901 = _zz_11902;
  assign _zz_11902 = ($signed(_zz_11903) >>> _zz_1676);
  assign _zz_11903 = _zz_11904;
  assign _zz_11904 = ($signed(data_mid_34_real) + $signed(_zz_1673));
  assign _zz_11905 = _zz_11906;
  assign _zz_11906 = ($signed(_zz_11907) >>> _zz_1676);
  assign _zz_11907 = _zz_11908;
  assign _zz_11908 = ($signed(data_mid_34_imag) + $signed(_zz_1674));
  assign _zz_11909 = ($signed(twiddle_factor_table_98_real) * $signed(data_mid_99_real));
  assign _zz_11910 = ($signed(twiddle_factor_table_98_imag) * $signed(data_mid_99_imag));
  assign _zz_11911 = fixTo_838_dout;
  assign _zz_11912 = ($signed(twiddle_factor_table_98_real) * $signed(data_mid_99_imag));
  assign _zz_11913 = ($signed(twiddle_factor_table_98_imag) * $signed(data_mid_99_real));
  assign _zz_11914 = fixTo_839_dout;
  assign _zz_11915 = _zz_11916;
  assign _zz_11916 = ($signed(_zz_11917) >>> _zz_1679);
  assign _zz_11917 = _zz_11918;
  assign _zz_11918 = ($signed(data_mid_35_real) - $signed(_zz_1677));
  assign _zz_11919 = _zz_11920;
  assign _zz_11920 = ($signed(_zz_11921) >>> _zz_1679);
  assign _zz_11921 = _zz_11922;
  assign _zz_11922 = ($signed(data_mid_35_imag) - $signed(_zz_1678));
  assign _zz_11923 = _zz_11924;
  assign _zz_11924 = ($signed(_zz_11925) >>> _zz_1680);
  assign _zz_11925 = _zz_11926;
  assign _zz_11926 = ($signed(data_mid_35_real) + $signed(_zz_1677));
  assign _zz_11927 = _zz_11928;
  assign _zz_11928 = ($signed(_zz_11929) >>> _zz_1680);
  assign _zz_11929 = _zz_11930;
  assign _zz_11930 = ($signed(data_mid_35_imag) + $signed(_zz_1678));
  assign _zz_11931 = ($signed(twiddle_factor_table_99_real) * $signed(data_mid_100_real));
  assign _zz_11932 = ($signed(twiddle_factor_table_99_imag) * $signed(data_mid_100_imag));
  assign _zz_11933 = fixTo_840_dout;
  assign _zz_11934 = ($signed(twiddle_factor_table_99_real) * $signed(data_mid_100_imag));
  assign _zz_11935 = ($signed(twiddle_factor_table_99_imag) * $signed(data_mid_100_real));
  assign _zz_11936 = fixTo_841_dout;
  assign _zz_11937 = _zz_11938;
  assign _zz_11938 = ($signed(_zz_11939) >>> _zz_1683);
  assign _zz_11939 = _zz_11940;
  assign _zz_11940 = ($signed(data_mid_36_real) - $signed(_zz_1681));
  assign _zz_11941 = _zz_11942;
  assign _zz_11942 = ($signed(_zz_11943) >>> _zz_1683);
  assign _zz_11943 = _zz_11944;
  assign _zz_11944 = ($signed(data_mid_36_imag) - $signed(_zz_1682));
  assign _zz_11945 = _zz_11946;
  assign _zz_11946 = ($signed(_zz_11947) >>> _zz_1684);
  assign _zz_11947 = _zz_11948;
  assign _zz_11948 = ($signed(data_mid_36_real) + $signed(_zz_1681));
  assign _zz_11949 = _zz_11950;
  assign _zz_11950 = ($signed(_zz_11951) >>> _zz_1684);
  assign _zz_11951 = _zz_11952;
  assign _zz_11952 = ($signed(data_mid_36_imag) + $signed(_zz_1682));
  assign _zz_11953 = ($signed(twiddle_factor_table_100_real) * $signed(data_mid_101_real));
  assign _zz_11954 = ($signed(twiddle_factor_table_100_imag) * $signed(data_mid_101_imag));
  assign _zz_11955 = fixTo_842_dout;
  assign _zz_11956 = ($signed(twiddle_factor_table_100_real) * $signed(data_mid_101_imag));
  assign _zz_11957 = ($signed(twiddle_factor_table_100_imag) * $signed(data_mid_101_real));
  assign _zz_11958 = fixTo_843_dout;
  assign _zz_11959 = _zz_11960;
  assign _zz_11960 = ($signed(_zz_11961) >>> _zz_1687);
  assign _zz_11961 = _zz_11962;
  assign _zz_11962 = ($signed(data_mid_37_real) - $signed(_zz_1685));
  assign _zz_11963 = _zz_11964;
  assign _zz_11964 = ($signed(_zz_11965) >>> _zz_1687);
  assign _zz_11965 = _zz_11966;
  assign _zz_11966 = ($signed(data_mid_37_imag) - $signed(_zz_1686));
  assign _zz_11967 = _zz_11968;
  assign _zz_11968 = ($signed(_zz_11969) >>> _zz_1688);
  assign _zz_11969 = _zz_11970;
  assign _zz_11970 = ($signed(data_mid_37_real) + $signed(_zz_1685));
  assign _zz_11971 = _zz_11972;
  assign _zz_11972 = ($signed(_zz_11973) >>> _zz_1688);
  assign _zz_11973 = _zz_11974;
  assign _zz_11974 = ($signed(data_mid_37_imag) + $signed(_zz_1686));
  assign _zz_11975 = ($signed(twiddle_factor_table_101_real) * $signed(data_mid_102_real));
  assign _zz_11976 = ($signed(twiddle_factor_table_101_imag) * $signed(data_mid_102_imag));
  assign _zz_11977 = fixTo_844_dout;
  assign _zz_11978 = ($signed(twiddle_factor_table_101_real) * $signed(data_mid_102_imag));
  assign _zz_11979 = ($signed(twiddle_factor_table_101_imag) * $signed(data_mid_102_real));
  assign _zz_11980 = fixTo_845_dout;
  assign _zz_11981 = _zz_11982;
  assign _zz_11982 = ($signed(_zz_11983) >>> _zz_1691);
  assign _zz_11983 = _zz_11984;
  assign _zz_11984 = ($signed(data_mid_38_real) - $signed(_zz_1689));
  assign _zz_11985 = _zz_11986;
  assign _zz_11986 = ($signed(_zz_11987) >>> _zz_1691);
  assign _zz_11987 = _zz_11988;
  assign _zz_11988 = ($signed(data_mid_38_imag) - $signed(_zz_1690));
  assign _zz_11989 = _zz_11990;
  assign _zz_11990 = ($signed(_zz_11991) >>> _zz_1692);
  assign _zz_11991 = _zz_11992;
  assign _zz_11992 = ($signed(data_mid_38_real) + $signed(_zz_1689));
  assign _zz_11993 = _zz_11994;
  assign _zz_11994 = ($signed(_zz_11995) >>> _zz_1692);
  assign _zz_11995 = _zz_11996;
  assign _zz_11996 = ($signed(data_mid_38_imag) + $signed(_zz_1690));
  assign _zz_11997 = ($signed(twiddle_factor_table_102_real) * $signed(data_mid_103_real));
  assign _zz_11998 = ($signed(twiddle_factor_table_102_imag) * $signed(data_mid_103_imag));
  assign _zz_11999 = fixTo_846_dout;
  assign _zz_12000 = ($signed(twiddle_factor_table_102_real) * $signed(data_mid_103_imag));
  assign _zz_12001 = ($signed(twiddle_factor_table_102_imag) * $signed(data_mid_103_real));
  assign _zz_12002 = fixTo_847_dout;
  assign _zz_12003 = _zz_12004;
  assign _zz_12004 = ($signed(_zz_12005) >>> _zz_1695);
  assign _zz_12005 = _zz_12006;
  assign _zz_12006 = ($signed(data_mid_39_real) - $signed(_zz_1693));
  assign _zz_12007 = _zz_12008;
  assign _zz_12008 = ($signed(_zz_12009) >>> _zz_1695);
  assign _zz_12009 = _zz_12010;
  assign _zz_12010 = ($signed(data_mid_39_imag) - $signed(_zz_1694));
  assign _zz_12011 = _zz_12012;
  assign _zz_12012 = ($signed(_zz_12013) >>> _zz_1696);
  assign _zz_12013 = _zz_12014;
  assign _zz_12014 = ($signed(data_mid_39_real) + $signed(_zz_1693));
  assign _zz_12015 = _zz_12016;
  assign _zz_12016 = ($signed(_zz_12017) >>> _zz_1696);
  assign _zz_12017 = _zz_12018;
  assign _zz_12018 = ($signed(data_mid_39_imag) + $signed(_zz_1694));
  assign _zz_12019 = ($signed(twiddle_factor_table_103_real) * $signed(data_mid_104_real));
  assign _zz_12020 = ($signed(twiddle_factor_table_103_imag) * $signed(data_mid_104_imag));
  assign _zz_12021 = fixTo_848_dout;
  assign _zz_12022 = ($signed(twiddle_factor_table_103_real) * $signed(data_mid_104_imag));
  assign _zz_12023 = ($signed(twiddle_factor_table_103_imag) * $signed(data_mid_104_real));
  assign _zz_12024 = fixTo_849_dout;
  assign _zz_12025 = _zz_12026;
  assign _zz_12026 = ($signed(_zz_12027) >>> _zz_1699);
  assign _zz_12027 = _zz_12028;
  assign _zz_12028 = ($signed(data_mid_40_real) - $signed(_zz_1697));
  assign _zz_12029 = _zz_12030;
  assign _zz_12030 = ($signed(_zz_12031) >>> _zz_1699);
  assign _zz_12031 = _zz_12032;
  assign _zz_12032 = ($signed(data_mid_40_imag) - $signed(_zz_1698));
  assign _zz_12033 = _zz_12034;
  assign _zz_12034 = ($signed(_zz_12035) >>> _zz_1700);
  assign _zz_12035 = _zz_12036;
  assign _zz_12036 = ($signed(data_mid_40_real) + $signed(_zz_1697));
  assign _zz_12037 = _zz_12038;
  assign _zz_12038 = ($signed(_zz_12039) >>> _zz_1700);
  assign _zz_12039 = _zz_12040;
  assign _zz_12040 = ($signed(data_mid_40_imag) + $signed(_zz_1698));
  assign _zz_12041 = ($signed(twiddle_factor_table_104_real) * $signed(data_mid_105_real));
  assign _zz_12042 = ($signed(twiddle_factor_table_104_imag) * $signed(data_mid_105_imag));
  assign _zz_12043 = fixTo_850_dout;
  assign _zz_12044 = ($signed(twiddle_factor_table_104_real) * $signed(data_mid_105_imag));
  assign _zz_12045 = ($signed(twiddle_factor_table_104_imag) * $signed(data_mid_105_real));
  assign _zz_12046 = fixTo_851_dout;
  assign _zz_12047 = _zz_12048;
  assign _zz_12048 = ($signed(_zz_12049) >>> _zz_1703);
  assign _zz_12049 = _zz_12050;
  assign _zz_12050 = ($signed(data_mid_41_real) - $signed(_zz_1701));
  assign _zz_12051 = _zz_12052;
  assign _zz_12052 = ($signed(_zz_12053) >>> _zz_1703);
  assign _zz_12053 = _zz_12054;
  assign _zz_12054 = ($signed(data_mid_41_imag) - $signed(_zz_1702));
  assign _zz_12055 = _zz_12056;
  assign _zz_12056 = ($signed(_zz_12057) >>> _zz_1704);
  assign _zz_12057 = _zz_12058;
  assign _zz_12058 = ($signed(data_mid_41_real) + $signed(_zz_1701));
  assign _zz_12059 = _zz_12060;
  assign _zz_12060 = ($signed(_zz_12061) >>> _zz_1704);
  assign _zz_12061 = _zz_12062;
  assign _zz_12062 = ($signed(data_mid_41_imag) + $signed(_zz_1702));
  assign _zz_12063 = ($signed(twiddle_factor_table_105_real) * $signed(data_mid_106_real));
  assign _zz_12064 = ($signed(twiddle_factor_table_105_imag) * $signed(data_mid_106_imag));
  assign _zz_12065 = fixTo_852_dout;
  assign _zz_12066 = ($signed(twiddle_factor_table_105_real) * $signed(data_mid_106_imag));
  assign _zz_12067 = ($signed(twiddle_factor_table_105_imag) * $signed(data_mid_106_real));
  assign _zz_12068 = fixTo_853_dout;
  assign _zz_12069 = _zz_12070;
  assign _zz_12070 = ($signed(_zz_12071) >>> _zz_1707);
  assign _zz_12071 = _zz_12072;
  assign _zz_12072 = ($signed(data_mid_42_real) - $signed(_zz_1705));
  assign _zz_12073 = _zz_12074;
  assign _zz_12074 = ($signed(_zz_12075) >>> _zz_1707);
  assign _zz_12075 = _zz_12076;
  assign _zz_12076 = ($signed(data_mid_42_imag) - $signed(_zz_1706));
  assign _zz_12077 = _zz_12078;
  assign _zz_12078 = ($signed(_zz_12079) >>> _zz_1708);
  assign _zz_12079 = _zz_12080;
  assign _zz_12080 = ($signed(data_mid_42_real) + $signed(_zz_1705));
  assign _zz_12081 = _zz_12082;
  assign _zz_12082 = ($signed(_zz_12083) >>> _zz_1708);
  assign _zz_12083 = _zz_12084;
  assign _zz_12084 = ($signed(data_mid_42_imag) + $signed(_zz_1706));
  assign _zz_12085 = ($signed(twiddle_factor_table_106_real) * $signed(data_mid_107_real));
  assign _zz_12086 = ($signed(twiddle_factor_table_106_imag) * $signed(data_mid_107_imag));
  assign _zz_12087 = fixTo_854_dout;
  assign _zz_12088 = ($signed(twiddle_factor_table_106_real) * $signed(data_mid_107_imag));
  assign _zz_12089 = ($signed(twiddle_factor_table_106_imag) * $signed(data_mid_107_real));
  assign _zz_12090 = fixTo_855_dout;
  assign _zz_12091 = _zz_12092;
  assign _zz_12092 = ($signed(_zz_12093) >>> _zz_1711);
  assign _zz_12093 = _zz_12094;
  assign _zz_12094 = ($signed(data_mid_43_real) - $signed(_zz_1709));
  assign _zz_12095 = _zz_12096;
  assign _zz_12096 = ($signed(_zz_12097) >>> _zz_1711);
  assign _zz_12097 = _zz_12098;
  assign _zz_12098 = ($signed(data_mid_43_imag) - $signed(_zz_1710));
  assign _zz_12099 = _zz_12100;
  assign _zz_12100 = ($signed(_zz_12101) >>> _zz_1712);
  assign _zz_12101 = _zz_12102;
  assign _zz_12102 = ($signed(data_mid_43_real) + $signed(_zz_1709));
  assign _zz_12103 = _zz_12104;
  assign _zz_12104 = ($signed(_zz_12105) >>> _zz_1712);
  assign _zz_12105 = _zz_12106;
  assign _zz_12106 = ($signed(data_mid_43_imag) + $signed(_zz_1710));
  assign _zz_12107 = ($signed(twiddle_factor_table_107_real) * $signed(data_mid_108_real));
  assign _zz_12108 = ($signed(twiddle_factor_table_107_imag) * $signed(data_mid_108_imag));
  assign _zz_12109 = fixTo_856_dout;
  assign _zz_12110 = ($signed(twiddle_factor_table_107_real) * $signed(data_mid_108_imag));
  assign _zz_12111 = ($signed(twiddle_factor_table_107_imag) * $signed(data_mid_108_real));
  assign _zz_12112 = fixTo_857_dout;
  assign _zz_12113 = _zz_12114;
  assign _zz_12114 = ($signed(_zz_12115) >>> _zz_1715);
  assign _zz_12115 = _zz_12116;
  assign _zz_12116 = ($signed(data_mid_44_real) - $signed(_zz_1713));
  assign _zz_12117 = _zz_12118;
  assign _zz_12118 = ($signed(_zz_12119) >>> _zz_1715);
  assign _zz_12119 = _zz_12120;
  assign _zz_12120 = ($signed(data_mid_44_imag) - $signed(_zz_1714));
  assign _zz_12121 = _zz_12122;
  assign _zz_12122 = ($signed(_zz_12123) >>> _zz_1716);
  assign _zz_12123 = _zz_12124;
  assign _zz_12124 = ($signed(data_mid_44_real) + $signed(_zz_1713));
  assign _zz_12125 = _zz_12126;
  assign _zz_12126 = ($signed(_zz_12127) >>> _zz_1716);
  assign _zz_12127 = _zz_12128;
  assign _zz_12128 = ($signed(data_mid_44_imag) + $signed(_zz_1714));
  assign _zz_12129 = ($signed(twiddle_factor_table_108_real) * $signed(data_mid_109_real));
  assign _zz_12130 = ($signed(twiddle_factor_table_108_imag) * $signed(data_mid_109_imag));
  assign _zz_12131 = fixTo_858_dout;
  assign _zz_12132 = ($signed(twiddle_factor_table_108_real) * $signed(data_mid_109_imag));
  assign _zz_12133 = ($signed(twiddle_factor_table_108_imag) * $signed(data_mid_109_real));
  assign _zz_12134 = fixTo_859_dout;
  assign _zz_12135 = _zz_12136;
  assign _zz_12136 = ($signed(_zz_12137) >>> _zz_1719);
  assign _zz_12137 = _zz_12138;
  assign _zz_12138 = ($signed(data_mid_45_real) - $signed(_zz_1717));
  assign _zz_12139 = _zz_12140;
  assign _zz_12140 = ($signed(_zz_12141) >>> _zz_1719);
  assign _zz_12141 = _zz_12142;
  assign _zz_12142 = ($signed(data_mid_45_imag) - $signed(_zz_1718));
  assign _zz_12143 = _zz_12144;
  assign _zz_12144 = ($signed(_zz_12145) >>> _zz_1720);
  assign _zz_12145 = _zz_12146;
  assign _zz_12146 = ($signed(data_mid_45_real) + $signed(_zz_1717));
  assign _zz_12147 = _zz_12148;
  assign _zz_12148 = ($signed(_zz_12149) >>> _zz_1720);
  assign _zz_12149 = _zz_12150;
  assign _zz_12150 = ($signed(data_mid_45_imag) + $signed(_zz_1718));
  assign _zz_12151 = ($signed(twiddle_factor_table_109_real) * $signed(data_mid_110_real));
  assign _zz_12152 = ($signed(twiddle_factor_table_109_imag) * $signed(data_mid_110_imag));
  assign _zz_12153 = fixTo_860_dout;
  assign _zz_12154 = ($signed(twiddle_factor_table_109_real) * $signed(data_mid_110_imag));
  assign _zz_12155 = ($signed(twiddle_factor_table_109_imag) * $signed(data_mid_110_real));
  assign _zz_12156 = fixTo_861_dout;
  assign _zz_12157 = _zz_12158;
  assign _zz_12158 = ($signed(_zz_12159) >>> _zz_1723);
  assign _zz_12159 = _zz_12160;
  assign _zz_12160 = ($signed(data_mid_46_real) - $signed(_zz_1721));
  assign _zz_12161 = _zz_12162;
  assign _zz_12162 = ($signed(_zz_12163) >>> _zz_1723);
  assign _zz_12163 = _zz_12164;
  assign _zz_12164 = ($signed(data_mid_46_imag) - $signed(_zz_1722));
  assign _zz_12165 = _zz_12166;
  assign _zz_12166 = ($signed(_zz_12167) >>> _zz_1724);
  assign _zz_12167 = _zz_12168;
  assign _zz_12168 = ($signed(data_mid_46_real) + $signed(_zz_1721));
  assign _zz_12169 = _zz_12170;
  assign _zz_12170 = ($signed(_zz_12171) >>> _zz_1724);
  assign _zz_12171 = _zz_12172;
  assign _zz_12172 = ($signed(data_mid_46_imag) + $signed(_zz_1722));
  assign _zz_12173 = ($signed(twiddle_factor_table_110_real) * $signed(data_mid_111_real));
  assign _zz_12174 = ($signed(twiddle_factor_table_110_imag) * $signed(data_mid_111_imag));
  assign _zz_12175 = fixTo_862_dout;
  assign _zz_12176 = ($signed(twiddle_factor_table_110_real) * $signed(data_mid_111_imag));
  assign _zz_12177 = ($signed(twiddle_factor_table_110_imag) * $signed(data_mid_111_real));
  assign _zz_12178 = fixTo_863_dout;
  assign _zz_12179 = _zz_12180;
  assign _zz_12180 = ($signed(_zz_12181) >>> _zz_1727);
  assign _zz_12181 = _zz_12182;
  assign _zz_12182 = ($signed(data_mid_47_real) - $signed(_zz_1725));
  assign _zz_12183 = _zz_12184;
  assign _zz_12184 = ($signed(_zz_12185) >>> _zz_1727);
  assign _zz_12185 = _zz_12186;
  assign _zz_12186 = ($signed(data_mid_47_imag) - $signed(_zz_1726));
  assign _zz_12187 = _zz_12188;
  assign _zz_12188 = ($signed(_zz_12189) >>> _zz_1728);
  assign _zz_12189 = _zz_12190;
  assign _zz_12190 = ($signed(data_mid_47_real) + $signed(_zz_1725));
  assign _zz_12191 = _zz_12192;
  assign _zz_12192 = ($signed(_zz_12193) >>> _zz_1728);
  assign _zz_12193 = _zz_12194;
  assign _zz_12194 = ($signed(data_mid_47_imag) + $signed(_zz_1726));
  assign _zz_12195 = ($signed(twiddle_factor_table_111_real) * $signed(data_mid_112_real));
  assign _zz_12196 = ($signed(twiddle_factor_table_111_imag) * $signed(data_mid_112_imag));
  assign _zz_12197 = fixTo_864_dout;
  assign _zz_12198 = ($signed(twiddle_factor_table_111_real) * $signed(data_mid_112_imag));
  assign _zz_12199 = ($signed(twiddle_factor_table_111_imag) * $signed(data_mid_112_real));
  assign _zz_12200 = fixTo_865_dout;
  assign _zz_12201 = _zz_12202;
  assign _zz_12202 = ($signed(_zz_12203) >>> _zz_1731);
  assign _zz_12203 = _zz_12204;
  assign _zz_12204 = ($signed(data_mid_48_real) - $signed(_zz_1729));
  assign _zz_12205 = _zz_12206;
  assign _zz_12206 = ($signed(_zz_12207) >>> _zz_1731);
  assign _zz_12207 = _zz_12208;
  assign _zz_12208 = ($signed(data_mid_48_imag) - $signed(_zz_1730));
  assign _zz_12209 = _zz_12210;
  assign _zz_12210 = ($signed(_zz_12211) >>> _zz_1732);
  assign _zz_12211 = _zz_12212;
  assign _zz_12212 = ($signed(data_mid_48_real) + $signed(_zz_1729));
  assign _zz_12213 = _zz_12214;
  assign _zz_12214 = ($signed(_zz_12215) >>> _zz_1732);
  assign _zz_12215 = _zz_12216;
  assign _zz_12216 = ($signed(data_mid_48_imag) + $signed(_zz_1730));
  assign _zz_12217 = ($signed(twiddle_factor_table_112_real) * $signed(data_mid_113_real));
  assign _zz_12218 = ($signed(twiddle_factor_table_112_imag) * $signed(data_mid_113_imag));
  assign _zz_12219 = fixTo_866_dout;
  assign _zz_12220 = ($signed(twiddle_factor_table_112_real) * $signed(data_mid_113_imag));
  assign _zz_12221 = ($signed(twiddle_factor_table_112_imag) * $signed(data_mid_113_real));
  assign _zz_12222 = fixTo_867_dout;
  assign _zz_12223 = _zz_12224;
  assign _zz_12224 = ($signed(_zz_12225) >>> _zz_1735);
  assign _zz_12225 = _zz_12226;
  assign _zz_12226 = ($signed(data_mid_49_real) - $signed(_zz_1733));
  assign _zz_12227 = _zz_12228;
  assign _zz_12228 = ($signed(_zz_12229) >>> _zz_1735);
  assign _zz_12229 = _zz_12230;
  assign _zz_12230 = ($signed(data_mid_49_imag) - $signed(_zz_1734));
  assign _zz_12231 = _zz_12232;
  assign _zz_12232 = ($signed(_zz_12233) >>> _zz_1736);
  assign _zz_12233 = _zz_12234;
  assign _zz_12234 = ($signed(data_mid_49_real) + $signed(_zz_1733));
  assign _zz_12235 = _zz_12236;
  assign _zz_12236 = ($signed(_zz_12237) >>> _zz_1736);
  assign _zz_12237 = _zz_12238;
  assign _zz_12238 = ($signed(data_mid_49_imag) + $signed(_zz_1734));
  assign _zz_12239 = ($signed(twiddle_factor_table_113_real) * $signed(data_mid_114_real));
  assign _zz_12240 = ($signed(twiddle_factor_table_113_imag) * $signed(data_mid_114_imag));
  assign _zz_12241 = fixTo_868_dout;
  assign _zz_12242 = ($signed(twiddle_factor_table_113_real) * $signed(data_mid_114_imag));
  assign _zz_12243 = ($signed(twiddle_factor_table_113_imag) * $signed(data_mid_114_real));
  assign _zz_12244 = fixTo_869_dout;
  assign _zz_12245 = _zz_12246;
  assign _zz_12246 = ($signed(_zz_12247) >>> _zz_1739);
  assign _zz_12247 = _zz_12248;
  assign _zz_12248 = ($signed(data_mid_50_real) - $signed(_zz_1737));
  assign _zz_12249 = _zz_12250;
  assign _zz_12250 = ($signed(_zz_12251) >>> _zz_1739);
  assign _zz_12251 = _zz_12252;
  assign _zz_12252 = ($signed(data_mid_50_imag) - $signed(_zz_1738));
  assign _zz_12253 = _zz_12254;
  assign _zz_12254 = ($signed(_zz_12255) >>> _zz_1740);
  assign _zz_12255 = _zz_12256;
  assign _zz_12256 = ($signed(data_mid_50_real) + $signed(_zz_1737));
  assign _zz_12257 = _zz_12258;
  assign _zz_12258 = ($signed(_zz_12259) >>> _zz_1740);
  assign _zz_12259 = _zz_12260;
  assign _zz_12260 = ($signed(data_mid_50_imag) + $signed(_zz_1738));
  assign _zz_12261 = ($signed(twiddle_factor_table_114_real) * $signed(data_mid_115_real));
  assign _zz_12262 = ($signed(twiddle_factor_table_114_imag) * $signed(data_mid_115_imag));
  assign _zz_12263 = fixTo_870_dout;
  assign _zz_12264 = ($signed(twiddle_factor_table_114_real) * $signed(data_mid_115_imag));
  assign _zz_12265 = ($signed(twiddle_factor_table_114_imag) * $signed(data_mid_115_real));
  assign _zz_12266 = fixTo_871_dout;
  assign _zz_12267 = _zz_12268;
  assign _zz_12268 = ($signed(_zz_12269) >>> _zz_1743);
  assign _zz_12269 = _zz_12270;
  assign _zz_12270 = ($signed(data_mid_51_real) - $signed(_zz_1741));
  assign _zz_12271 = _zz_12272;
  assign _zz_12272 = ($signed(_zz_12273) >>> _zz_1743);
  assign _zz_12273 = _zz_12274;
  assign _zz_12274 = ($signed(data_mid_51_imag) - $signed(_zz_1742));
  assign _zz_12275 = _zz_12276;
  assign _zz_12276 = ($signed(_zz_12277) >>> _zz_1744);
  assign _zz_12277 = _zz_12278;
  assign _zz_12278 = ($signed(data_mid_51_real) + $signed(_zz_1741));
  assign _zz_12279 = _zz_12280;
  assign _zz_12280 = ($signed(_zz_12281) >>> _zz_1744);
  assign _zz_12281 = _zz_12282;
  assign _zz_12282 = ($signed(data_mid_51_imag) + $signed(_zz_1742));
  assign _zz_12283 = ($signed(twiddle_factor_table_115_real) * $signed(data_mid_116_real));
  assign _zz_12284 = ($signed(twiddle_factor_table_115_imag) * $signed(data_mid_116_imag));
  assign _zz_12285 = fixTo_872_dout;
  assign _zz_12286 = ($signed(twiddle_factor_table_115_real) * $signed(data_mid_116_imag));
  assign _zz_12287 = ($signed(twiddle_factor_table_115_imag) * $signed(data_mid_116_real));
  assign _zz_12288 = fixTo_873_dout;
  assign _zz_12289 = _zz_12290;
  assign _zz_12290 = ($signed(_zz_12291) >>> _zz_1747);
  assign _zz_12291 = _zz_12292;
  assign _zz_12292 = ($signed(data_mid_52_real) - $signed(_zz_1745));
  assign _zz_12293 = _zz_12294;
  assign _zz_12294 = ($signed(_zz_12295) >>> _zz_1747);
  assign _zz_12295 = _zz_12296;
  assign _zz_12296 = ($signed(data_mid_52_imag) - $signed(_zz_1746));
  assign _zz_12297 = _zz_12298;
  assign _zz_12298 = ($signed(_zz_12299) >>> _zz_1748);
  assign _zz_12299 = _zz_12300;
  assign _zz_12300 = ($signed(data_mid_52_real) + $signed(_zz_1745));
  assign _zz_12301 = _zz_12302;
  assign _zz_12302 = ($signed(_zz_12303) >>> _zz_1748);
  assign _zz_12303 = _zz_12304;
  assign _zz_12304 = ($signed(data_mid_52_imag) + $signed(_zz_1746));
  assign _zz_12305 = ($signed(twiddle_factor_table_116_real) * $signed(data_mid_117_real));
  assign _zz_12306 = ($signed(twiddle_factor_table_116_imag) * $signed(data_mid_117_imag));
  assign _zz_12307 = fixTo_874_dout;
  assign _zz_12308 = ($signed(twiddle_factor_table_116_real) * $signed(data_mid_117_imag));
  assign _zz_12309 = ($signed(twiddle_factor_table_116_imag) * $signed(data_mid_117_real));
  assign _zz_12310 = fixTo_875_dout;
  assign _zz_12311 = _zz_12312;
  assign _zz_12312 = ($signed(_zz_12313) >>> _zz_1751);
  assign _zz_12313 = _zz_12314;
  assign _zz_12314 = ($signed(data_mid_53_real) - $signed(_zz_1749));
  assign _zz_12315 = _zz_12316;
  assign _zz_12316 = ($signed(_zz_12317) >>> _zz_1751);
  assign _zz_12317 = _zz_12318;
  assign _zz_12318 = ($signed(data_mid_53_imag) - $signed(_zz_1750));
  assign _zz_12319 = _zz_12320;
  assign _zz_12320 = ($signed(_zz_12321) >>> _zz_1752);
  assign _zz_12321 = _zz_12322;
  assign _zz_12322 = ($signed(data_mid_53_real) + $signed(_zz_1749));
  assign _zz_12323 = _zz_12324;
  assign _zz_12324 = ($signed(_zz_12325) >>> _zz_1752);
  assign _zz_12325 = _zz_12326;
  assign _zz_12326 = ($signed(data_mid_53_imag) + $signed(_zz_1750));
  assign _zz_12327 = ($signed(twiddle_factor_table_117_real) * $signed(data_mid_118_real));
  assign _zz_12328 = ($signed(twiddle_factor_table_117_imag) * $signed(data_mid_118_imag));
  assign _zz_12329 = fixTo_876_dout;
  assign _zz_12330 = ($signed(twiddle_factor_table_117_real) * $signed(data_mid_118_imag));
  assign _zz_12331 = ($signed(twiddle_factor_table_117_imag) * $signed(data_mid_118_real));
  assign _zz_12332 = fixTo_877_dout;
  assign _zz_12333 = _zz_12334;
  assign _zz_12334 = ($signed(_zz_12335) >>> _zz_1755);
  assign _zz_12335 = _zz_12336;
  assign _zz_12336 = ($signed(data_mid_54_real) - $signed(_zz_1753));
  assign _zz_12337 = _zz_12338;
  assign _zz_12338 = ($signed(_zz_12339) >>> _zz_1755);
  assign _zz_12339 = _zz_12340;
  assign _zz_12340 = ($signed(data_mid_54_imag) - $signed(_zz_1754));
  assign _zz_12341 = _zz_12342;
  assign _zz_12342 = ($signed(_zz_12343) >>> _zz_1756);
  assign _zz_12343 = _zz_12344;
  assign _zz_12344 = ($signed(data_mid_54_real) + $signed(_zz_1753));
  assign _zz_12345 = _zz_12346;
  assign _zz_12346 = ($signed(_zz_12347) >>> _zz_1756);
  assign _zz_12347 = _zz_12348;
  assign _zz_12348 = ($signed(data_mid_54_imag) + $signed(_zz_1754));
  assign _zz_12349 = ($signed(twiddle_factor_table_118_real) * $signed(data_mid_119_real));
  assign _zz_12350 = ($signed(twiddle_factor_table_118_imag) * $signed(data_mid_119_imag));
  assign _zz_12351 = fixTo_878_dout;
  assign _zz_12352 = ($signed(twiddle_factor_table_118_real) * $signed(data_mid_119_imag));
  assign _zz_12353 = ($signed(twiddle_factor_table_118_imag) * $signed(data_mid_119_real));
  assign _zz_12354 = fixTo_879_dout;
  assign _zz_12355 = _zz_12356;
  assign _zz_12356 = ($signed(_zz_12357) >>> _zz_1759);
  assign _zz_12357 = _zz_12358;
  assign _zz_12358 = ($signed(data_mid_55_real) - $signed(_zz_1757));
  assign _zz_12359 = _zz_12360;
  assign _zz_12360 = ($signed(_zz_12361) >>> _zz_1759);
  assign _zz_12361 = _zz_12362;
  assign _zz_12362 = ($signed(data_mid_55_imag) - $signed(_zz_1758));
  assign _zz_12363 = _zz_12364;
  assign _zz_12364 = ($signed(_zz_12365) >>> _zz_1760);
  assign _zz_12365 = _zz_12366;
  assign _zz_12366 = ($signed(data_mid_55_real) + $signed(_zz_1757));
  assign _zz_12367 = _zz_12368;
  assign _zz_12368 = ($signed(_zz_12369) >>> _zz_1760);
  assign _zz_12369 = _zz_12370;
  assign _zz_12370 = ($signed(data_mid_55_imag) + $signed(_zz_1758));
  assign _zz_12371 = ($signed(twiddle_factor_table_119_real) * $signed(data_mid_120_real));
  assign _zz_12372 = ($signed(twiddle_factor_table_119_imag) * $signed(data_mid_120_imag));
  assign _zz_12373 = fixTo_880_dout;
  assign _zz_12374 = ($signed(twiddle_factor_table_119_real) * $signed(data_mid_120_imag));
  assign _zz_12375 = ($signed(twiddle_factor_table_119_imag) * $signed(data_mid_120_real));
  assign _zz_12376 = fixTo_881_dout;
  assign _zz_12377 = _zz_12378;
  assign _zz_12378 = ($signed(_zz_12379) >>> _zz_1763);
  assign _zz_12379 = _zz_12380;
  assign _zz_12380 = ($signed(data_mid_56_real) - $signed(_zz_1761));
  assign _zz_12381 = _zz_12382;
  assign _zz_12382 = ($signed(_zz_12383) >>> _zz_1763);
  assign _zz_12383 = _zz_12384;
  assign _zz_12384 = ($signed(data_mid_56_imag) - $signed(_zz_1762));
  assign _zz_12385 = _zz_12386;
  assign _zz_12386 = ($signed(_zz_12387) >>> _zz_1764);
  assign _zz_12387 = _zz_12388;
  assign _zz_12388 = ($signed(data_mid_56_real) + $signed(_zz_1761));
  assign _zz_12389 = _zz_12390;
  assign _zz_12390 = ($signed(_zz_12391) >>> _zz_1764);
  assign _zz_12391 = _zz_12392;
  assign _zz_12392 = ($signed(data_mid_56_imag) + $signed(_zz_1762));
  assign _zz_12393 = ($signed(twiddle_factor_table_120_real) * $signed(data_mid_121_real));
  assign _zz_12394 = ($signed(twiddle_factor_table_120_imag) * $signed(data_mid_121_imag));
  assign _zz_12395 = fixTo_882_dout;
  assign _zz_12396 = ($signed(twiddle_factor_table_120_real) * $signed(data_mid_121_imag));
  assign _zz_12397 = ($signed(twiddle_factor_table_120_imag) * $signed(data_mid_121_real));
  assign _zz_12398 = fixTo_883_dout;
  assign _zz_12399 = _zz_12400;
  assign _zz_12400 = ($signed(_zz_12401) >>> _zz_1767);
  assign _zz_12401 = _zz_12402;
  assign _zz_12402 = ($signed(data_mid_57_real) - $signed(_zz_1765));
  assign _zz_12403 = _zz_12404;
  assign _zz_12404 = ($signed(_zz_12405) >>> _zz_1767);
  assign _zz_12405 = _zz_12406;
  assign _zz_12406 = ($signed(data_mid_57_imag) - $signed(_zz_1766));
  assign _zz_12407 = _zz_12408;
  assign _zz_12408 = ($signed(_zz_12409) >>> _zz_1768);
  assign _zz_12409 = _zz_12410;
  assign _zz_12410 = ($signed(data_mid_57_real) + $signed(_zz_1765));
  assign _zz_12411 = _zz_12412;
  assign _zz_12412 = ($signed(_zz_12413) >>> _zz_1768);
  assign _zz_12413 = _zz_12414;
  assign _zz_12414 = ($signed(data_mid_57_imag) + $signed(_zz_1766));
  assign _zz_12415 = ($signed(twiddle_factor_table_121_real) * $signed(data_mid_122_real));
  assign _zz_12416 = ($signed(twiddle_factor_table_121_imag) * $signed(data_mid_122_imag));
  assign _zz_12417 = fixTo_884_dout;
  assign _zz_12418 = ($signed(twiddle_factor_table_121_real) * $signed(data_mid_122_imag));
  assign _zz_12419 = ($signed(twiddle_factor_table_121_imag) * $signed(data_mid_122_real));
  assign _zz_12420 = fixTo_885_dout;
  assign _zz_12421 = _zz_12422;
  assign _zz_12422 = ($signed(_zz_12423) >>> _zz_1771);
  assign _zz_12423 = _zz_12424;
  assign _zz_12424 = ($signed(data_mid_58_real) - $signed(_zz_1769));
  assign _zz_12425 = _zz_12426;
  assign _zz_12426 = ($signed(_zz_12427) >>> _zz_1771);
  assign _zz_12427 = _zz_12428;
  assign _zz_12428 = ($signed(data_mid_58_imag) - $signed(_zz_1770));
  assign _zz_12429 = _zz_12430;
  assign _zz_12430 = ($signed(_zz_12431) >>> _zz_1772);
  assign _zz_12431 = _zz_12432;
  assign _zz_12432 = ($signed(data_mid_58_real) + $signed(_zz_1769));
  assign _zz_12433 = _zz_12434;
  assign _zz_12434 = ($signed(_zz_12435) >>> _zz_1772);
  assign _zz_12435 = _zz_12436;
  assign _zz_12436 = ($signed(data_mid_58_imag) + $signed(_zz_1770));
  assign _zz_12437 = ($signed(twiddle_factor_table_122_real) * $signed(data_mid_123_real));
  assign _zz_12438 = ($signed(twiddle_factor_table_122_imag) * $signed(data_mid_123_imag));
  assign _zz_12439 = fixTo_886_dout;
  assign _zz_12440 = ($signed(twiddle_factor_table_122_real) * $signed(data_mid_123_imag));
  assign _zz_12441 = ($signed(twiddle_factor_table_122_imag) * $signed(data_mid_123_real));
  assign _zz_12442 = fixTo_887_dout;
  assign _zz_12443 = _zz_12444;
  assign _zz_12444 = ($signed(_zz_12445) >>> _zz_1775);
  assign _zz_12445 = _zz_12446;
  assign _zz_12446 = ($signed(data_mid_59_real) - $signed(_zz_1773));
  assign _zz_12447 = _zz_12448;
  assign _zz_12448 = ($signed(_zz_12449) >>> _zz_1775);
  assign _zz_12449 = _zz_12450;
  assign _zz_12450 = ($signed(data_mid_59_imag) - $signed(_zz_1774));
  assign _zz_12451 = _zz_12452;
  assign _zz_12452 = ($signed(_zz_12453) >>> _zz_1776);
  assign _zz_12453 = _zz_12454;
  assign _zz_12454 = ($signed(data_mid_59_real) + $signed(_zz_1773));
  assign _zz_12455 = _zz_12456;
  assign _zz_12456 = ($signed(_zz_12457) >>> _zz_1776);
  assign _zz_12457 = _zz_12458;
  assign _zz_12458 = ($signed(data_mid_59_imag) + $signed(_zz_1774));
  assign _zz_12459 = ($signed(twiddle_factor_table_123_real) * $signed(data_mid_124_real));
  assign _zz_12460 = ($signed(twiddle_factor_table_123_imag) * $signed(data_mid_124_imag));
  assign _zz_12461 = fixTo_888_dout;
  assign _zz_12462 = ($signed(twiddle_factor_table_123_real) * $signed(data_mid_124_imag));
  assign _zz_12463 = ($signed(twiddle_factor_table_123_imag) * $signed(data_mid_124_real));
  assign _zz_12464 = fixTo_889_dout;
  assign _zz_12465 = _zz_12466;
  assign _zz_12466 = ($signed(_zz_12467) >>> _zz_1779);
  assign _zz_12467 = _zz_12468;
  assign _zz_12468 = ($signed(data_mid_60_real) - $signed(_zz_1777));
  assign _zz_12469 = _zz_12470;
  assign _zz_12470 = ($signed(_zz_12471) >>> _zz_1779);
  assign _zz_12471 = _zz_12472;
  assign _zz_12472 = ($signed(data_mid_60_imag) - $signed(_zz_1778));
  assign _zz_12473 = _zz_12474;
  assign _zz_12474 = ($signed(_zz_12475) >>> _zz_1780);
  assign _zz_12475 = _zz_12476;
  assign _zz_12476 = ($signed(data_mid_60_real) + $signed(_zz_1777));
  assign _zz_12477 = _zz_12478;
  assign _zz_12478 = ($signed(_zz_12479) >>> _zz_1780);
  assign _zz_12479 = _zz_12480;
  assign _zz_12480 = ($signed(data_mid_60_imag) + $signed(_zz_1778));
  assign _zz_12481 = ($signed(twiddle_factor_table_124_real) * $signed(data_mid_125_real));
  assign _zz_12482 = ($signed(twiddle_factor_table_124_imag) * $signed(data_mid_125_imag));
  assign _zz_12483 = fixTo_890_dout;
  assign _zz_12484 = ($signed(twiddle_factor_table_124_real) * $signed(data_mid_125_imag));
  assign _zz_12485 = ($signed(twiddle_factor_table_124_imag) * $signed(data_mid_125_real));
  assign _zz_12486 = fixTo_891_dout;
  assign _zz_12487 = _zz_12488;
  assign _zz_12488 = ($signed(_zz_12489) >>> _zz_1783);
  assign _zz_12489 = _zz_12490;
  assign _zz_12490 = ($signed(data_mid_61_real) - $signed(_zz_1781));
  assign _zz_12491 = _zz_12492;
  assign _zz_12492 = ($signed(_zz_12493) >>> _zz_1783);
  assign _zz_12493 = _zz_12494;
  assign _zz_12494 = ($signed(data_mid_61_imag) - $signed(_zz_1782));
  assign _zz_12495 = _zz_12496;
  assign _zz_12496 = ($signed(_zz_12497) >>> _zz_1784);
  assign _zz_12497 = _zz_12498;
  assign _zz_12498 = ($signed(data_mid_61_real) + $signed(_zz_1781));
  assign _zz_12499 = _zz_12500;
  assign _zz_12500 = ($signed(_zz_12501) >>> _zz_1784);
  assign _zz_12501 = _zz_12502;
  assign _zz_12502 = ($signed(data_mid_61_imag) + $signed(_zz_1782));
  assign _zz_12503 = ($signed(twiddle_factor_table_125_real) * $signed(data_mid_126_real));
  assign _zz_12504 = ($signed(twiddle_factor_table_125_imag) * $signed(data_mid_126_imag));
  assign _zz_12505 = fixTo_892_dout;
  assign _zz_12506 = ($signed(twiddle_factor_table_125_real) * $signed(data_mid_126_imag));
  assign _zz_12507 = ($signed(twiddle_factor_table_125_imag) * $signed(data_mid_126_real));
  assign _zz_12508 = fixTo_893_dout;
  assign _zz_12509 = _zz_12510;
  assign _zz_12510 = ($signed(_zz_12511) >>> _zz_1787);
  assign _zz_12511 = _zz_12512;
  assign _zz_12512 = ($signed(data_mid_62_real) - $signed(_zz_1785));
  assign _zz_12513 = _zz_12514;
  assign _zz_12514 = ($signed(_zz_12515) >>> _zz_1787);
  assign _zz_12515 = _zz_12516;
  assign _zz_12516 = ($signed(data_mid_62_imag) - $signed(_zz_1786));
  assign _zz_12517 = _zz_12518;
  assign _zz_12518 = ($signed(_zz_12519) >>> _zz_1788);
  assign _zz_12519 = _zz_12520;
  assign _zz_12520 = ($signed(data_mid_62_real) + $signed(_zz_1785));
  assign _zz_12521 = _zz_12522;
  assign _zz_12522 = ($signed(_zz_12523) >>> _zz_1788);
  assign _zz_12523 = _zz_12524;
  assign _zz_12524 = ($signed(data_mid_62_imag) + $signed(_zz_1786));
  assign _zz_12525 = ($signed(twiddle_factor_table_126_real) * $signed(data_mid_127_real));
  assign _zz_12526 = ($signed(twiddle_factor_table_126_imag) * $signed(data_mid_127_imag));
  assign _zz_12527 = fixTo_894_dout;
  assign _zz_12528 = ($signed(twiddle_factor_table_126_real) * $signed(data_mid_127_imag));
  assign _zz_12529 = ($signed(twiddle_factor_table_126_imag) * $signed(data_mid_127_real));
  assign _zz_12530 = fixTo_895_dout;
  assign _zz_12531 = _zz_12532;
  assign _zz_12532 = ($signed(_zz_12533) >>> _zz_1791);
  assign _zz_12533 = _zz_12534;
  assign _zz_12534 = ($signed(data_mid_63_real) - $signed(_zz_1789));
  assign _zz_12535 = _zz_12536;
  assign _zz_12536 = ($signed(_zz_12537) >>> _zz_1791);
  assign _zz_12537 = _zz_12538;
  assign _zz_12538 = ($signed(data_mid_63_imag) - $signed(_zz_1790));
  assign _zz_12539 = _zz_12540;
  assign _zz_12540 = ($signed(_zz_12541) >>> _zz_1792);
  assign _zz_12541 = _zz_12542;
  assign _zz_12542 = ($signed(data_mid_63_real) + $signed(_zz_1789));
  assign _zz_12543 = _zz_12544;
  assign _zz_12544 = ($signed(_zz_12545) >>> _zz_1792);
  assign _zz_12545 = _zz_12546;
  assign _zz_12546 = ($signed(data_mid_63_imag) + $signed(_zz_1790));
  SInt32fixTo23_8_ROUNDTOINF fixTo (
    .din     (_zz_1793[31:0]    ), //i
    .dout    (fixTo_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1 (
    .din     (_zz_1794[31:0]      ), //i
    .dout    (fixTo_1_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2 (
    .din     (_zz_1795[31:0]      ), //i
    .dout    (fixTo_2_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_3 (
    .din     (_zz_1796[31:0]      ), //i
    .dout    (fixTo_3_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_4 (
    .din     (_zz_1797[31:0]      ), //i
    .dout    (fixTo_4_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_5 (
    .din     (_zz_1798[31:0]      ), //i
    .dout    (fixTo_5_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_6 (
    .din     (_zz_1799[31:0]      ), //i
    .dout    (fixTo_6_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_7 (
    .din     (_zz_1800[31:0]      ), //i
    .dout    (fixTo_7_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_8 (
    .din     (_zz_1801[31:0]      ), //i
    .dout    (fixTo_8_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_9 (
    .din     (_zz_1802[31:0]      ), //i
    .dout    (fixTo_9_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_10 (
    .din     (_zz_1803[31:0]       ), //i
    .dout    (fixTo_10_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_11 (
    .din     (_zz_1804[31:0]       ), //i
    .dout    (fixTo_11_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_12 (
    .din     (_zz_1805[31:0]       ), //i
    .dout    (fixTo_12_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_13 (
    .din     (_zz_1806[31:0]       ), //i
    .dout    (fixTo_13_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_14 (
    .din     (_zz_1807[31:0]       ), //i
    .dout    (fixTo_14_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_15 (
    .din     (_zz_1808[31:0]       ), //i
    .dout    (fixTo_15_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_16 (
    .din     (_zz_1809[31:0]       ), //i
    .dout    (fixTo_16_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_17 (
    .din     (_zz_1810[31:0]       ), //i
    .dout    (fixTo_17_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_18 (
    .din     (_zz_1811[31:0]       ), //i
    .dout    (fixTo_18_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_19 (
    .din     (_zz_1812[31:0]       ), //i
    .dout    (fixTo_19_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_20 (
    .din     (_zz_1813[31:0]       ), //i
    .dout    (fixTo_20_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_21 (
    .din     (_zz_1814[31:0]       ), //i
    .dout    (fixTo_21_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_22 (
    .din     (_zz_1815[31:0]       ), //i
    .dout    (fixTo_22_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_23 (
    .din     (_zz_1816[31:0]       ), //i
    .dout    (fixTo_23_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_24 (
    .din     (_zz_1817[31:0]       ), //i
    .dout    (fixTo_24_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_25 (
    .din     (_zz_1818[31:0]       ), //i
    .dout    (fixTo_25_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_26 (
    .din     (_zz_1819[31:0]       ), //i
    .dout    (fixTo_26_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_27 (
    .din     (_zz_1820[31:0]       ), //i
    .dout    (fixTo_27_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_28 (
    .din     (_zz_1821[31:0]       ), //i
    .dout    (fixTo_28_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_29 (
    .din     (_zz_1822[31:0]       ), //i
    .dout    (fixTo_29_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_30 (
    .din     (_zz_1823[31:0]       ), //i
    .dout    (fixTo_30_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_31 (
    .din     (_zz_1824[31:0]       ), //i
    .dout    (fixTo_31_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_32 (
    .din     (_zz_1825[31:0]       ), //i
    .dout    (fixTo_32_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_33 (
    .din     (_zz_1826[31:0]       ), //i
    .dout    (fixTo_33_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_34 (
    .din     (_zz_1827[31:0]       ), //i
    .dout    (fixTo_34_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_35 (
    .din     (_zz_1828[31:0]       ), //i
    .dout    (fixTo_35_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_36 (
    .din     (_zz_1829[31:0]       ), //i
    .dout    (fixTo_36_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_37 (
    .din     (_zz_1830[31:0]       ), //i
    .dout    (fixTo_37_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_38 (
    .din     (_zz_1831[31:0]       ), //i
    .dout    (fixTo_38_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_39 (
    .din     (_zz_1832[31:0]       ), //i
    .dout    (fixTo_39_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_40 (
    .din     (_zz_1833[31:0]       ), //i
    .dout    (fixTo_40_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_41 (
    .din     (_zz_1834[31:0]       ), //i
    .dout    (fixTo_41_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_42 (
    .din     (_zz_1835[31:0]       ), //i
    .dout    (fixTo_42_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_43 (
    .din     (_zz_1836[31:0]       ), //i
    .dout    (fixTo_43_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_44 (
    .din     (_zz_1837[31:0]       ), //i
    .dout    (fixTo_44_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_45 (
    .din     (_zz_1838[31:0]       ), //i
    .dout    (fixTo_45_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_46 (
    .din     (_zz_1839[31:0]       ), //i
    .dout    (fixTo_46_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_47 (
    .din     (_zz_1840[31:0]       ), //i
    .dout    (fixTo_47_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_48 (
    .din     (_zz_1841[31:0]       ), //i
    .dout    (fixTo_48_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_49 (
    .din     (_zz_1842[31:0]       ), //i
    .dout    (fixTo_49_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_50 (
    .din     (_zz_1843[31:0]       ), //i
    .dout    (fixTo_50_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_51 (
    .din     (_zz_1844[31:0]       ), //i
    .dout    (fixTo_51_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_52 (
    .din     (_zz_1845[31:0]       ), //i
    .dout    (fixTo_52_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_53 (
    .din     (_zz_1846[31:0]       ), //i
    .dout    (fixTo_53_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_54 (
    .din     (_zz_1847[31:0]       ), //i
    .dout    (fixTo_54_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_55 (
    .din     (_zz_1848[31:0]       ), //i
    .dout    (fixTo_55_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_56 (
    .din     (_zz_1849[31:0]       ), //i
    .dout    (fixTo_56_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_57 (
    .din     (_zz_1850[31:0]       ), //i
    .dout    (fixTo_57_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_58 (
    .din     (_zz_1851[31:0]       ), //i
    .dout    (fixTo_58_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_59 (
    .din     (_zz_1852[31:0]       ), //i
    .dout    (fixTo_59_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_60 (
    .din     (_zz_1853[31:0]       ), //i
    .dout    (fixTo_60_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_61 (
    .din     (_zz_1854[31:0]       ), //i
    .dout    (fixTo_61_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_62 (
    .din     (_zz_1855[31:0]       ), //i
    .dout    (fixTo_62_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_63 (
    .din     (_zz_1856[31:0]       ), //i
    .dout    (fixTo_63_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_64 (
    .din     (_zz_1857[31:0]       ), //i
    .dout    (fixTo_64_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_65 (
    .din     (_zz_1858[31:0]       ), //i
    .dout    (fixTo_65_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_66 (
    .din     (_zz_1859[31:0]       ), //i
    .dout    (fixTo_66_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_67 (
    .din     (_zz_1860[31:0]       ), //i
    .dout    (fixTo_67_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_68 (
    .din     (_zz_1861[31:0]       ), //i
    .dout    (fixTo_68_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_69 (
    .din     (_zz_1862[31:0]       ), //i
    .dout    (fixTo_69_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_70 (
    .din     (_zz_1863[31:0]       ), //i
    .dout    (fixTo_70_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_71 (
    .din     (_zz_1864[31:0]       ), //i
    .dout    (fixTo_71_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_72 (
    .din     (_zz_1865[31:0]       ), //i
    .dout    (fixTo_72_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_73 (
    .din     (_zz_1866[31:0]       ), //i
    .dout    (fixTo_73_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_74 (
    .din     (_zz_1867[31:0]       ), //i
    .dout    (fixTo_74_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_75 (
    .din     (_zz_1868[31:0]       ), //i
    .dout    (fixTo_75_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_76 (
    .din     (_zz_1869[31:0]       ), //i
    .dout    (fixTo_76_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_77 (
    .din     (_zz_1870[31:0]       ), //i
    .dout    (fixTo_77_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_78 (
    .din     (_zz_1871[31:0]       ), //i
    .dout    (fixTo_78_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_79 (
    .din     (_zz_1872[31:0]       ), //i
    .dout    (fixTo_79_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_80 (
    .din     (_zz_1873[31:0]       ), //i
    .dout    (fixTo_80_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_81 (
    .din     (_zz_1874[31:0]       ), //i
    .dout    (fixTo_81_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_82 (
    .din     (_zz_1875[31:0]       ), //i
    .dout    (fixTo_82_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_83 (
    .din     (_zz_1876[31:0]       ), //i
    .dout    (fixTo_83_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_84 (
    .din     (_zz_1877[31:0]       ), //i
    .dout    (fixTo_84_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_85 (
    .din     (_zz_1878[31:0]       ), //i
    .dout    (fixTo_85_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_86 (
    .din     (_zz_1879[31:0]       ), //i
    .dout    (fixTo_86_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_87 (
    .din     (_zz_1880[31:0]       ), //i
    .dout    (fixTo_87_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_88 (
    .din     (_zz_1881[31:0]       ), //i
    .dout    (fixTo_88_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_89 (
    .din     (_zz_1882[31:0]       ), //i
    .dout    (fixTo_89_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_90 (
    .din     (_zz_1883[31:0]       ), //i
    .dout    (fixTo_90_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_91 (
    .din     (_zz_1884[31:0]       ), //i
    .dout    (fixTo_91_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_92 (
    .din     (_zz_1885[31:0]       ), //i
    .dout    (fixTo_92_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_93 (
    .din     (_zz_1886[31:0]       ), //i
    .dout    (fixTo_93_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_94 (
    .din     (_zz_1887[31:0]       ), //i
    .dout    (fixTo_94_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_95 (
    .din     (_zz_1888[31:0]       ), //i
    .dout    (fixTo_95_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_96 (
    .din     (_zz_1889[31:0]       ), //i
    .dout    (fixTo_96_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_97 (
    .din     (_zz_1890[31:0]       ), //i
    .dout    (fixTo_97_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_98 (
    .din     (_zz_1891[31:0]       ), //i
    .dout    (fixTo_98_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_99 (
    .din     (_zz_1892[31:0]       ), //i
    .dout    (fixTo_99_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_100 (
    .din     (_zz_1893[31:0]        ), //i
    .dout    (fixTo_100_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_101 (
    .din     (_zz_1894[31:0]        ), //i
    .dout    (fixTo_101_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_102 (
    .din     (_zz_1895[31:0]        ), //i
    .dout    (fixTo_102_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_103 (
    .din     (_zz_1896[31:0]        ), //i
    .dout    (fixTo_103_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_104 (
    .din     (_zz_1897[31:0]        ), //i
    .dout    (fixTo_104_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_105 (
    .din     (_zz_1898[31:0]        ), //i
    .dout    (fixTo_105_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_106 (
    .din     (_zz_1899[31:0]        ), //i
    .dout    (fixTo_106_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_107 (
    .din     (_zz_1900[31:0]        ), //i
    .dout    (fixTo_107_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_108 (
    .din     (_zz_1901[31:0]        ), //i
    .dout    (fixTo_108_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_109 (
    .din     (_zz_1902[31:0]        ), //i
    .dout    (fixTo_109_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_110 (
    .din     (_zz_1903[31:0]        ), //i
    .dout    (fixTo_110_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_111 (
    .din     (_zz_1904[31:0]        ), //i
    .dout    (fixTo_111_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_112 (
    .din     (_zz_1905[31:0]        ), //i
    .dout    (fixTo_112_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_113 (
    .din     (_zz_1906[31:0]        ), //i
    .dout    (fixTo_113_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_114 (
    .din     (_zz_1907[31:0]        ), //i
    .dout    (fixTo_114_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_115 (
    .din     (_zz_1908[31:0]        ), //i
    .dout    (fixTo_115_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_116 (
    .din     (_zz_1909[31:0]        ), //i
    .dout    (fixTo_116_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_117 (
    .din     (_zz_1910[31:0]        ), //i
    .dout    (fixTo_117_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_118 (
    .din     (_zz_1911[31:0]        ), //i
    .dout    (fixTo_118_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_119 (
    .din     (_zz_1912[31:0]        ), //i
    .dout    (fixTo_119_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_120 (
    .din     (_zz_1913[31:0]        ), //i
    .dout    (fixTo_120_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_121 (
    .din     (_zz_1914[31:0]        ), //i
    .dout    (fixTo_121_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_122 (
    .din     (_zz_1915[31:0]        ), //i
    .dout    (fixTo_122_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_123 (
    .din     (_zz_1916[31:0]        ), //i
    .dout    (fixTo_123_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_124 (
    .din     (_zz_1917[31:0]        ), //i
    .dout    (fixTo_124_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_125 (
    .din     (_zz_1918[31:0]        ), //i
    .dout    (fixTo_125_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_126 (
    .din     (_zz_1919[31:0]        ), //i
    .dout    (fixTo_126_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_127 (
    .din     (_zz_1920[31:0]        ), //i
    .dout    (fixTo_127_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_128 (
    .din     (_zz_1921[31:0]        ), //i
    .dout    (fixTo_128_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_129 (
    .din     (_zz_1922[31:0]        ), //i
    .dout    (fixTo_129_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_130 (
    .din     (_zz_1923[31:0]        ), //i
    .dout    (fixTo_130_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_131 (
    .din     (_zz_1924[31:0]        ), //i
    .dout    (fixTo_131_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_132 (
    .din     (_zz_1925[31:0]        ), //i
    .dout    (fixTo_132_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_133 (
    .din     (_zz_1926[31:0]        ), //i
    .dout    (fixTo_133_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_134 (
    .din     (_zz_1927[31:0]        ), //i
    .dout    (fixTo_134_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_135 (
    .din     (_zz_1928[31:0]        ), //i
    .dout    (fixTo_135_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_136 (
    .din     (_zz_1929[31:0]        ), //i
    .dout    (fixTo_136_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_137 (
    .din     (_zz_1930[31:0]        ), //i
    .dout    (fixTo_137_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_138 (
    .din     (_zz_1931[31:0]        ), //i
    .dout    (fixTo_138_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_139 (
    .din     (_zz_1932[31:0]        ), //i
    .dout    (fixTo_139_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_140 (
    .din     (_zz_1933[31:0]        ), //i
    .dout    (fixTo_140_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_141 (
    .din     (_zz_1934[31:0]        ), //i
    .dout    (fixTo_141_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_142 (
    .din     (_zz_1935[31:0]        ), //i
    .dout    (fixTo_142_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_143 (
    .din     (_zz_1936[31:0]        ), //i
    .dout    (fixTo_143_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_144 (
    .din     (_zz_1937[31:0]        ), //i
    .dout    (fixTo_144_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_145 (
    .din     (_zz_1938[31:0]        ), //i
    .dout    (fixTo_145_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_146 (
    .din     (_zz_1939[31:0]        ), //i
    .dout    (fixTo_146_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_147 (
    .din     (_zz_1940[31:0]        ), //i
    .dout    (fixTo_147_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_148 (
    .din     (_zz_1941[31:0]        ), //i
    .dout    (fixTo_148_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_149 (
    .din     (_zz_1942[31:0]        ), //i
    .dout    (fixTo_149_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_150 (
    .din     (_zz_1943[31:0]        ), //i
    .dout    (fixTo_150_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_151 (
    .din     (_zz_1944[31:0]        ), //i
    .dout    (fixTo_151_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_152 (
    .din     (_zz_1945[31:0]        ), //i
    .dout    (fixTo_152_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_153 (
    .din     (_zz_1946[31:0]        ), //i
    .dout    (fixTo_153_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_154 (
    .din     (_zz_1947[31:0]        ), //i
    .dout    (fixTo_154_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_155 (
    .din     (_zz_1948[31:0]        ), //i
    .dout    (fixTo_155_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_156 (
    .din     (_zz_1949[31:0]        ), //i
    .dout    (fixTo_156_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_157 (
    .din     (_zz_1950[31:0]        ), //i
    .dout    (fixTo_157_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_158 (
    .din     (_zz_1951[31:0]        ), //i
    .dout    (fixTo_158_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_159 (
    .din     (_zz_1952[31:0]        ), //i
    .dout    (fixTo_159_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_160 (
    .din     (_zz_1953[31:0]        ), //i
    .dout    (fixTo_160_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_161 (
    .din     (_zz_1954[31:0]        ), //i
    .dout    (fixTo_161_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_162 (
    .din     (_zz_1955[31:0]        ), //i
    .dout    (fixTo_162_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_163 (
    .din     (_zz_1956[31:0]        ), //i
    .dout    (fixTo_163_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_164 (
    .din     (_zz_1957[31:0]        ), //i
    .dout    (fixTo_164_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_165 (
    .din     (_zz_1958[31:0]        ), //i
    .dout    (fixTo_165_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_166 (
    .din     (_zz_1959[31:0]        ), //i
    .dout    (fixTo_166_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_167 (
    .din     (_zz_1960[31:0]        ), //i
    .dout    (fixTo_167_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_168 (
    .din     (_zz_1961[31:0]        ), //i
    .dout    (fixTo_168_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_169 (
    .din     (_zz_1962[31:0]        ), //i
    .dout    (fixTo_169_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_170 (
    .din     (_zz_1963[31:0]        ), //i
    .dout    (fixTo_170_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_171 (
    .din     (_zz_1964[31:0]        ), //i
    .dout    (fixTo_171_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_172 (
    .din     (_zz_1965[31:0]        ), //i
    .dout    (fixTo_172_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_173 (
    .din     (_zz_1966[31:0]        ), //i
    .dout    (fixTo_173_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_174 (
    .din     (_zz_1967[31:0]        ), //i
    .dout    (fixTo_174_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_175 (
    .din     (_zz_1968[31:0]        ), //i
    .dout    (fixTo_175_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_176 (
    .din     (_zz_1969[31:0]        ), //i
    .dout    (fixTo_176_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_177 (
    .din     (_zz_1970[31:0]        ), //i
    .dout    (fixTo_177_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_178 (
    .din     (_zz_1971[31:0]        ), //i
    .dout    (fixTo_178_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_179 (
    .din     (_zz_1972[31:0]        ), //i
    .dout    (fixTo_179_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_180 (
    .din     (_zz_1973[31:0]        ), //i
    .dout    (fixTo_180_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_181 (
    .din     (_zz_1974[31:0]        ), //i
    .dout    (fixTo_181_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_182 (
    .din     (_zz_1975[31:0]        ), //i
    .dout    (fixTo_182_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_183 (
    .din     (_zz_1976[31:0]        ), //i
    .dout    (fixTo_183_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_184 (
    .din     (_zz_1977[31:0]        ), //i
    .dout    (fixTo_184_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_185 (
    .din     (_zz_1978[31:0]        ), //i
    .dout    (fixTo_185_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_186 (
    .din     (_zz_1979[31:0]        ), //i
    .dout    (fixTo_186_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_187 (
    .din     (_zz_1980[31:0]        ), //i
    .dout    (fixTo_187_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_188 (
    .din     (_zz_1981[31:0]        ), //i
    .dout    (fixTo_188_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_189 (
    .din     (_zz_1982[31:0]        ), //i
    .dout    (fixTo_189_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_190 (
    .din     (_zz_1983[31:0]        ), //i
    .dout    (fixTo_190_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_191 (
    .din     (_zz_1984[31:0]        ), //i
    .dout    (fixTo_191_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_192 (
    .din     (_zz_1985[31:0]        ), //i
    .dout    (fixTo_192_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_193 (
    .din     (_zz_1986[31:0]        ), //i
    .dout    (fixTo_193_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_194 (
    .din     (_zz_1987[31:0]        ), //i
    .dout    (fixTo_194_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_195 (
    .din     (_zz_1988[31:0]        ), //i
    .dout    (fixTo_195_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_196 (
    .din     (_zz_1989[31:0]        ), //i
    .dout    (fixTo_196_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_197 (
    .din     (_zz_1990[31:0]        ), //i
    .dout    (fixTo_197_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_198 (
    .din     (_zz_1991[31:0]        ), //i
    .dout    (fixTo_198_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_199 (
    .din     (_zz_1992[31:0]        ), //i
    .dout    (fixTo_199_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_200 (
    .din     (_zz_1993[31:0]        ), //i
    .dout    (fixTo_200_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_201 (
    .din     (_zz_1994[31:0]        ), //i
    .dout    (fixTo_201_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_202 (
    .din     (_zz_1995[31:0]        ), //i
    .dout    (fixTo_202_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_203 (
    .din     (_zz_1996[31:0]        ), //i
    .dout    (fixTo_203_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_204 (
    .din     (_zz_1997[31:0]        ), //i
    .dout    (fixTo_204_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_205 (
    .din     (_zz_1998[31:0]        ), //i
    .dout    (fixTo_205_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_206 (
    .din     (_zz_1999[31:0]        ), //i
    .dout    (fixTo_206_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_207 (
    .din     (_zz_2000[31:0]        ), //i
    .dout    (fixTo_207_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_208 (
    .din     (_zz_2001[31:0]        ), //i
    .dout    (fixTo_208_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_209 (
    .din     (_zz_2002[31:0]        ), //i
    .dout    (fixTo_209_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_210 (
    .din     (_zz_2003[31:0]        ), //i
    .dout    (fixTo_210_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_211 (
    .din     (_zz_2004[31:0]        ), //i
    .dout    (fixTo_211_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_212 (
    .din     (_zz_2005[31:0]        ), //i
    .dout    (fixTo_212_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_213 (
    .din     (_zz_2006[31:0]        ), //i
    .dout    (fixTo_213_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_214 (
    .din     (_zz_2007[31:0]        ), //i
    .dout    (fixTo_214_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_215 (
    .din     (_zz_2008[31:0]        ), //i
    .dout    (fixTo_215_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_216 (
    .din     (_zz_2009[31:0]        ), //i
    .dout    (fixTo_216_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_217 (
    .din     (_zz_2010[31:0]        ), //i
    .dout    (fixTo_217_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_218 (
    .din     (_zz_2011[31:0]        ), //i
    .dout    (fixTo_218_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_219 (
    .din     (_zz_2012[31:0]        ), //i
    .dout    (fixTo_219_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_220 (
    .din     (_zz_2013[31:0]        ), //i
    .dout    (fixTo_220_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_221 (
    .din     (_zz_2014[31:0]        ), //i
    .dout    (fixTo_221_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_222 (
    .din     (_zz_2015[31:0]        ), //i
    .dout    (fixTo_222_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_223 (
    .din     (_zz_2016[31:0]        ), //i
    .dout    (fixTo_223_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_224 (
    .din     (_zz_2017[31:0]        ), //i
    .dout    (fixTo_224_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_225 (
    .din     (_zz_2018[31:0]        ), //i
    .dout    (fixTo_225_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_226 (
    .din     (_zz_2019[31:0]        ), //i
    .dout    (fixTo_226_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_227 (
    .din     (_zz_2020[31:0]        ), //i
    .dout    (fixTo_227_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_228 (
    .din     (_zz_2021[31:0]        ), //i
    .dout    (fixTo_228_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_229 (
    .din     (_zz_2022[31:0]        ), //i
    .dout    (fixTo_229_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_230 (
    .din     (_zz_2023[31:0]        ), //i
    .dout    (fixTo_230_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_231 (
    .din     (_zz_2024[31:0]        ), //i
    .dout    (fixTo_231_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_232 (
    .din     (_zz_2025[31:0]        ), //i
    .dout    (fixTo_232_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_233 (
    .din     (_zz_2026[31:0]        ), //i
    .dout    (fixTo_233_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_234 (
    .din     (_zz_2027[31:0]        ), //i
    .dout    (fixTo_234_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_235 (
    .din     (_zz_2028[31:0]        ), //i
    .dout    (fixTo_235_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_236 (
    .din     (_zz_2029[31:0]        ), //i
    .dout    (fixTo_236_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_237 (
    .din     (_zz_2030[31:0]        ), //i
    .dout    (fixTo_237_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_238 (
    .din     (_zz_2031[31:0]        ), //i
    .dout    (fixTo_238_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_239 (
    .din     (_zz_2032[31:0]        ), //i
    .dout    (fixTo_239_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_240 (
    .din     (_zz_2033[31:0]        ), //i
    .dout    (fixTo_240_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_241 (
    .din     (_zz_2034[31:0]        ), //i
    .dout    (fixTo_241_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_242 (
    .din     (_zz_2035[31:0]        ), //i
    .dout    (fixTo_242_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_243 (
    .din     (_zz_2036[31:0]        ), //i
    .dout    (fixTo_243_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_244 (
    .din     (_zz_2037[31:0]        ), //i
    .dout    (fixTo_244_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_245 (
    .din     (_zz_2038[31:0]        ), //i
    .dout    (fixTo_245_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_246 (
    .din     (_zz_2039[31:0]        ), //i
    .dout    (fixTo_246_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_247 (
    .din     (_zz_2040[31:0]        ), //i
    .dout    (fixTo_247_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_248 (
    .din     (_zz_2041[31:0]        ), //i
    .dout    (fixTo_248_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_249 (
    .din     (_zz_2042[31:0]        ), //i
    .dout    (fixTo_249_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_250 (
    .din     (_zz_2043[31:0]        ), //i
    .dout    (fixTo_250_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_251 (
    .din     (_zz_2044[31:0]        ), //i
    .dout    (fixTo_251_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_252 (
    .din     (_zz_2045[31:0]        ), //i
    .dout    (fixTo_252_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_253 (
    .din     (_zz_2046[31:0]        ), //i
    .dout    (fixTo_253_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_254 (
    .din     (_zz_2047[31:0]        ), //i
    .dout    (fixTo_254_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_255 (
    .din     (_zz_2048[31:0]        ), //i
    .dout    (fixTo_255_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_256 (
    .din     (_zz_2049[31:0]        ), //i
    .dout    (fixTo_256_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_257 (
    .din     (_zz_2050[31:0]        ), //i
    .dout    (fixTo_257_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_258 (
    .din     (_zz_2051[31:0]        ), //i
    .dout    (fixTo_258_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_259 (
    .din     (_zz_2052[31:0]        ), //i
    .dout    (fixTo_259_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_260 (
    .din     (_zz_2053[31:0]        ), //i
    .dout    (fixTo_260_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_261 (
    .din     (_zz_2054[31:0]        ), //i
    .dout    (fixTo_261_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_262 (
    .din     (_zz_2055[31:0]        ), //i
    .dout    (fixTo_262_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_263 (
    .din     (_zz_2056[31:0]        ), //i
    .dout    (fixTo_263_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_264 (
    .din     (_zz_2057[31:0]        ), //i
    .dout    (fixTo_264_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_265 (
    .din     (_zz_2058[31:0]        ), //i
    .dout    (fixTo_265_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_266 (
    .din     (_zz_2059[31:0]        ), //i
    .dout    (fixTo_266_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_267 (
    .din     (_zz_2060[31:0]        ), //i
    .dout    (fixTo_267_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_268 (
    .din     (_zz_2061[31:0]        ), //i
    .dout    (fixTo_268_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_269 (
    .din     (_zz_2062[31:0]        ), //i
    .dout    (fixTo_269_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_270 (
    .din     (_zz_2063[31:0]        ), //i
    .dout    (fixTo_270_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_271 (
    .din     (_zz_2064[31:0]        ), //i
    .dout    (fixTo_271_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_272 (
    .din     (_zz_2065[31:0]        ), //i
    .dout    (fixTo_272_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_273 (
    .din     (_zz_2066[31:0]        ), //i
    .dout    (fixTo_273_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_274 (
    .din     (_zz_2067[31:0]        ), //i
    .dout    (fixTo_274_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_275 (
    .din     (_zz_2068[31:0]        ), //i
    .dout    (fixTo_275_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_276 (
    .din     (_zz_2069[31:0]        ), //i
    .dout    (fixTo_276_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_277 (
    .din     (_zz_2070[31:0]        ), //i
    .dout    (fixTo_277_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_278 (
    .din     (_zz_2071[31:0]        ), //i
    .dout    (fixTo_278_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_279 (
    .din     (_zz_2072[31:0]        ), //i
    .dout    (fixTo_279_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_280 (
    .din     (_zz_2073[31:0]        ), //i
    .dout    (fixTo_280_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_281 (
    .din     (_zz_2074[31:0]        ), //i
    .dout    (fixTo_281_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_282 (
    .din     (_zz_2075[31:0]        ), //i
    .dout    (fixTo_282_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_283 (
    .din     (_zz_2076[31:0]        ), //i
    .dout    (fixTo_283_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_284 (
    .din     (_zz_2077[31:0]        ), //i
    .dout    (fixTo_284_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_285 (
    .din     (_zz_2078[31:0]        ), //i
    .dout    (fixTo_285_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_286 (
    .din     (_zz_2079[31:0]        ), //i
    .dout    (fixTo_286_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_287 (
    .din     (_zz_2080[31:0]        ), //i
    .dout    (fixTo_287_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_288 (
    .din     (_zz_2081[31:0]        ), //i
    .dout    (fixTo_288_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_289 (
    .din     (_zz_2082[31:0]        ), //i
    .dout    (fixTo_289_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_290 (
    .din     (_zz_2083[31:0]        ), //i
    .dout    (fixTo_290_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_291 (
    .din     (_zz_2084[31:0]        ), //i
    .dout    (fixTo_291_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_292 (
    .din     (_zz_2085[31:0]        ), //i
    .dout    (fixTo_292_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_293 (
    .din     (_zz_2086[31:0]        ), //i
    .dout    (fixTo_293_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_294 (
    .din     (_zz_2087[31:0]        ), //i
    .dout    (fixTo_294_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_295 (
    .din     (_zz_2088[31:0]        ), //i
    .dout    (fixTo_295_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_296 (
    .din     (_zz_2089[31:0]        ), //i
    .dout    (fixTo_296_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_297 (
    .din     (_zz_2090[31:0]        ), //i
    .dout    (fixTo_297_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_298 (
    .din     (_zz_2091[31:0]        ), //i
    .dout    (fixTo_298_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_299 (
    .din     (_zz_2092[31:0]        ), //i
    .dout    (fixTo_299_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_300 (
    .din     (_zz_2093[31:0]        ), //i
    .dout    (fixTo_300_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_301 (
    .din     (_zz_2094[31:0]        ), //i
    .dout    (fixTo_301_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_302 (
    .din     (_zz_2095[31:0]        ), //i
    .dout    (fixTo_302_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_303 (
    .din     (_zz_2096[31:0]        ), //i
    .dout    (fixTo_303_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_304 (
    .din     (_zz_2097[31:0]        ), //i
    .dout    (fixTo_304_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_305 (
    .din     (_zz_2098[31:0]        ), //i
    .dout    (fixTo_305_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_306 (
    .din     (_zz_2099[31:0]        ), //i
    .dout    (fixTo_306_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_307 (
    .din     (_zz_2100[31:0]        ), //i
    .dout    (fixTo_307_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_308 (
    .din     (_zz_2101[31:0]        ), //i
    .dout    (fixTo_308_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_309 (
    .din     (_zz_2102[31:0]        ), //i
    .dout    (fixTo_309_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_310 (
    .din     (_zz_2103[31:0]        ), //i
    .dout    (fixTo_310_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_311 (
    .din     (_zz_2104[31:0]        ), //i
    .dout    (fixTo_311_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_312 (
    .din     (_zz_2105[31:0]        ), //i
    .dout    (fixTo_312_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_313 (
    .din     (_zz_2106[31:0]        ), //i
    .dout    (fixTo_313_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_314 (
    .din     (_zz_2107[31:0]        ), //i
    .dout    (fixTo_314_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_315 (
    .din     (_zz_2108[31:0]        ), //i
    .dout    (fixTo_315_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_316 (
    .din     (_zz_2109[31:0]        ), //i
    .dout    (fixTo_316_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_317 (
    .din     (_zz_2110[31:0]        ), //i
    .dout    (fixTo_317_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_318 (
    .din     (_zz_2111[31:0]        ), //i
    .dout    (fixTo_318_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_319 (
    .din     (_zz_2112[31:0]        ), //i
    .dout    (fixTo_319_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_320 (
    .din     (_zz_2113[31:0]        ), //i
    .dout    (fixTo_320_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_321 (
    .din     (_zz_2114[31:0]        ), //i
    .dout    (fixTo_321_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_322 (
    .din     (_zz_2115[31:0]        ), //i
    .dout    (fixTo_322_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_323 (
    .din     (_zz_2116[31:0]        ), //i
    .dout    (fixTo_323_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_324 (
    .din     (_zz_2117[31:0]        ), //i
    .dout    (fixTo_324_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_325 (
    .din     (_zz_2118[31:0]        ), //i
    .dout    (fixTo_325_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_326 (
    .din     (_zz_2119[31:0]        ), //i
    .dout    (fixTo_326_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_327 (
    .din     (_zz_2120[31:0]        ), //i
    .dout    (fixTo_327_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_328 (
    .din     (_zz_2121[31:0]        ), //i
    .dout    (fixTo_328_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_329 (
    .din     (_zz_2122[31:0]        ), //i
    .dout    (fixTo_329_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_330 (
    .din     (_zz_2123[31:0]        ), //i
    .dout    (fixTo_330_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_331 (
    .din     (_zz_2124[31:0]        ), //i
    .dout    (fixTo_331_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_332 (
    .din     (_zz_2125[31:0]        ), //i
    .dout    (fixTo_332_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_333 (
    .din     (_zz_2126[31:0]        ), //i
    .dout    (fixTo_333_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_334 (
    .din     (_zz_2127[31:0]        ), //i
    .dout    (fixTo_334_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_335 (
    .din     (_zz_2128[31:0]        ), //i
    .dout    (fixTo_335_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_336 (
    .din     (_zz_2129[31:0]        ), //i
    .dout    (fixTo_336_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_337 (
    .din     (_zz_2130[31:0]        ), //i
    .dout    (fixTo_337_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_338 (
    .din     (_zz_2131[31:0]        ), //i
    .dout    (fixTo_338_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_339 (
    .din     (_zz_2132[31:0]        ), //i
    .dout    (fixTo_339_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_340 (
    .din     (_zz_2133[31:0]        ), //i
    .dout    (fixTo_340_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_341 (
    .din     (_zz_2134[31:0]        ), //i
    .dout    (fixTo_341_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_342 (
    .din     (_zz_2135[31:0]        ), //i
    .dout    (fixTo_342_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_343 (
    .din     (_zz_2136[31:0]        ), //i
    .dout    (fixTo_343_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_344 (
    .din     (_zz_2137[31:0]        ), //i
    .dout    (fixTo_344_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_345 (
    .din     (_zz_2138[31:0]        ), //i
    .dout    (fixTo_345_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_346 (
    .din     (_zz_2139[31:0]        ), //i
    .dout    (fixTo_346_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_347 (
    .din     (_zz_2140[31:0]        ), //i
    .dout    (fixTo_347_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_348 (
    .din     (_zz_2141[31:0]        ), //i
    .dout    (fixTo_348_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_349 (
    .din     (_zz_2142[31:0]        ), //i
    .dout    (fixTo_349_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_350 (
    .din     (_zz_2143[31:0]        ), //i
    .dout    (fixTo_350_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_351 (
    .din     (_zz_2144[31:0]        ), //i
    .dout    (fixTo_351_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_352 (
    .din     (_zz_2145[31:0]        ), //i
    .dout    (fixTo_352_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_353 (
    .din     (_zz_2146[31:0]        ), //i
    .dout    (fixTo_353_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_354 (
    .din     (_zz_2147[31:0]        ), //i
    .dout    (fixTo_354_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_355 (
    .din     (_zz_2148[31:0]        ), //i
    .dout    (fixTo_355_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_356 (
    .din     (_zz_2149[31:0]        ), //i
    .dout    (fixTo_356_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_357 (
    .din     (_zz_2150[31:0]        ), //i
    .dout    (fixTo_357_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_358 (
    .din     (_zz_2151[31:0]        ), //i
    .dout    (fixTo_358_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_359 (
    .din     (_zz_2152[31:0]        ), //i
    .dout    (fixTo_359_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_360 (
    .din     (_zz_2153[31:0]        ), //i
    .dout    (fixTo_360_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_361 (
    .din     (_zz_2154[31:0]        ), //i
    .dout    (fixTo_361_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_362 (
    .din     (_zz_2155[31:0]        ), //i
    .dout    (fixTo_362_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_363 (
    .din     (_zz_2156[31:0]        ), //i
    .dout    (fixTo_363_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_364 (
    .din     (_zz_2157[31:0]        ), //i
    .dout    (fixTo_364_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_365 (
    .din     (_zz_2158[31:0]        ), //i
    .dout    (fixTo_365_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_366 (
    .din     (_zz_2159[31:0]        ), //i
    .dout    (fixTo_366_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_367 (
    .din     (_zz_2160[31:0]        ), //i
    .dout    (fixTo_367_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_368 (
    .din     (_zz_2161[31:0]        ), //i
    .dout    (fixTo_368_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_369 (
    .din     (_zz_2162[31:0]        ), //i
    .dout    (fixTo_369_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_370 (
    .din     (_zz_2163[31:0]        ), //i
    .dout    (fixTo_370_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_371 (
    .din     (_zz_2164[31:0]        ), //i
    .dout    (fixTo_371_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_372 (
    .din     (_zz_2165[31:0]        ), //i
    .dout    (fixTo_372_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_373 (
    .din     (_zz_2166[31:0]        ), //i
    .dout    (fixTo_373_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_374 (
    .din     (_zz_2167[31:0]        ), //i
    .dout    (fixTo_374_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_375 (
    .din     (_zz_2168[31:0]        ), //i
    .dout    (fixTo_375_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_376 (
    .din     (_zz_2169[31:0]        ), //i
    .dout    (fixTo_376_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_377 (
    .din     (_zz_2170[31:0]        ), //i
    .dout    (fixTo_377_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_378 (
    .din     (_zz_2171[31:0]        ), //i
    .dout    (fixTo_378_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_379 (
    .din     (_zz_2172[31:0]        ), //i
    .dout    (fixTo_379_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_380 (
    .din     (_zz_2173[31:0]        ), //i
    .dout    (fixTo_380_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_381 (
    .din     (_zz_2174[31:0]        ), //i
    .dout    (fixTo_381_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_382 (
    .din     (_zz_2175[31:0]        ), //i
    .dout    (fixTo_382_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_383 (
    .din     (_zz_2176[31:0]        ), //i
    .dout    (fixTo_383_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_384 (
    .din     (_zz_2177[31:0]        ), //i
    .dout    (fixTo_384_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_385 (
    .din     (_zz_2178[31:0]        ), //i
    .dout    (fixTo_385_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_386 (
    .din     (_zz_2179[31:0]        ), //i
    .dout    (fixTo_386_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_387 (
    .din     (_zz_2180[31:0]        ), //i
    .dout    (fixTo_387_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_388 (
    .din     (_zz_2181[31:0]        ), //i
    .dout    (fixTo_388_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_389 (
    .din     (_zz_2182[31:0]        ), //i
    .dout    (fixTo_389_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_390 (
    .din     (_zz_2183[31:0]        ), //i
    .dout    (fixTo_390_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_391 (
    .din     (_zz_2184[31:0]        ), //i
    .dout    (fixTo_391_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_392 (
    .din     (_zz_2185[31:0]        ), //i
    .dout    (fixTo_392_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_393 (
    .din     (_zz_2186[31:0]        ), //i
    .dout    (fixTo_393_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_394 (
    .din     (_zz_2187[31:0]        ), //i
    .dout    (fixTo_394_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_395 (
    .din     (_zz_2188[31:0]        ), //i
    .dout    (fixTo_395_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_396 (
    .din     (_zz_2189[31:0]        ), //i
    .dout    (fixTo_396_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_397 (
    .din     (_zz_2190[31:0]        ), //i
    .dout    (fixTo_397_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_398 (
    .din     (_zz_2191[31:0]        ), //i
    .dout    (fixTo_398_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_399 (
    .din     (_zz_2192[31:0]        ), //i
    .dout    (fixTo_399_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_400 (
    .din     (_zz_2193[31:0]        ), //i
    .dout    (fixTo_400_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_401 (
    .din     (_zz_2194[31:0]        ), //i
    .dout    (fixTo_401_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_402 (
    .din     (_zz_2195[31:0]        ), //i
    .dout    (fixTo_402_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_403 (
    .din     (_zz_2196[31:0]        ), //i
    .dout    (fixTo_403_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_404 (
    .din     (_zz_2197[31:0]        ), //i
    .dout    (fixTo_404_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_405 (
    .din     (_zz_2198[31:0]        ), //i
    .dout    (fixTo_405_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_406 (
    .din     (_zz_2199[31:0]        ), //i
    .dout    (fixTo_406_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_407 (
    .din     (_zz_2200[31:0]        ), //i
    .dout    (fixTo_407_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_408 (
    .din     (_zz_2201[31:0]        ), //i
    .dout    (fixTo_408_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_409 (
    .din     (_zz_2202[31:0]        ), //i
    .dout    (fixTo_409_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_410 (
    .din     (_zz_2203[31:0]        ), //i
    .dout    (fixTo_410_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_411 (
    .din     (_zz_2204[31:0]        ), //i
    .dout    (fixTo_411_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_412 (
    .din     (_zz_2205[31:0]        ), //i
    .dout    (fixTo_412_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_413 (
    .din     (_zz_2206[31:0]        ), //i
    .dout    (fixTo_413_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_414 (
    .din     (_zz_2207[31:0]        ), //i
    .dout    (fixTo_414_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_415 (
    .din     (_zz_2208[31:0]        ), //i
    .dout    (fixTo_415_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_416 (
    .din     (_zz_2209[31:0]        ), //i
    .dout    (fixTo_416_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_417 (
    .din     (_zz_2210[31:0]        ), //i
    .dout    (fixTo_417_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_418 (
    .din     (_zz_2211[31:0]        ), //i
    .dout    (fixTo_418_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_419 (
    .din     (_zz_2212[31:0]        ), //i
    .dout    (fixTo_419_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_420 (
    .din     (_zz_2213[31:0]        ), //i
    .dout    (fixTo_420_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_421 (
    .din     (_zz_2214[31:0]        ), //i
    .dout    (fixTo_421_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_422 (
    .din     (_zz_2215[31:0]        ), //i
    .dout    (fixTo_422_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_423 (
    .din     (_zz_2216[31:0]        ), //i
    .dout    (fixTo_423_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_424 (
    .din     (_zz_2217[31:0]        ), //i
    .dout    (fixTo_424_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_425 (
    .din     (_zz_2218[31:0]        ), //i
    .dout    (fixTo_425_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_426 (
    .din     (_zz_2219[31:0]        ), //i
    .dout    (fixTo_426_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_427 (
    .din     (_zz_2220[31:0]        ), //i
    .dout    (fixTo_427_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_428 (
    .din     (_zz_2221[31:0]        ), //i
    .dout    (fixTo_428_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_429 (
    .din     (_zz_2222[31:0]        ), //i
    .dout    (fixTo_429_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_430 (
    .din     (_zz_2223[31:0]        ), //i
    .dout    (fixTo_430_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_431 (
    .din     (_zz_2224[31:0]        ), //i
    .dout    (fixTo_431_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_432 (
    .din     (_zz_2225[31:0]        ), //i
    .dout    (fixTo_432_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_433 (
    .din     (_zz_2226[31:0]        ), //i
    .dout    (fixTo_433_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_434 (
    .din     (_zz_2227[31:0]        ), //i
    .dout    (fixTo_434_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_435 (
    .din     (_zz_2228[31:0]        ), //i
    .dout    (fixTo_435_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_436 (
    .din     (_zz_2229[31:0]        ), //i
    .dout    (fixTo_436_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_437 (
    .din     (_zz_2230[31:0]        ), //i
    .dout    (fixTo_437_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_438 (
    .din     (_zz_2231[31:0]        ), //i
    .dout    (fixTo_438_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_439 (
    .din     (_zz_2232[31:0]        ), //i
    .dout    (fixTo_439_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_440 (
    .din     (_zz_2233[31:0]        ), //i
    .dout    (fixTo_440_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_441 (
    .din     (_zz_2234[31:0]        ), //i
    .dout    (fixTo_441_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_442 (
    .din     (_zz_2235[31:0]        ), //i
    .dout    (fixTo_442_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_443 (
    .din     (_zz_2236[31:0]        ), //i
    .dout    (fixTo_443_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_444 (
    .din     (_zz_2237[31:0]        ), //i
    .dout    (fixTo_444_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_445 (
    .din     (_zz_2238[31:0]        ), //i
    .dout    (fixTo_445_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_446 (
    .din     (_zz_2239[31:0]        ), //i
    .dout    (fixTo_446_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_447 (
    .din     (_zz_2240[31:0]        ), //i
    .dout    (fixTo_447_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_448 (
    .din     (_zz_2241[31:0]        ), //i
    .dout    (fixTo_448_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_449 (
    .din     (_zz_2242[31:0]        ), //i
    .dout    (fixTo_449_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_450 (
    .din     (_zz_2243[31:0]        ), //i
    .dout    (fixTo_450_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_451 (
    .din     (_zz_2244[31:0]        ), //i
    .dout    (fixTo_451_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_452 (
    .din     (_zz_2245[31:0]        ), //i
    .dout    (fixTo_452_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_453 (
    .din     (_zz_2246[31:0]        ), //i
    .dout    (fixTo_453_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_454 (
    .din     (_zz_2247[31:0]        ), //i
    .dout    (fixTo_454_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_455 (
    .din     (_zz_2248[31:0]        ), //i
    .dout    (fixTo_455_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_456 (
    .din     (_zz_2249[31:0]        ), //i
    .dout    (fixTo_456_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_457 (
    .din     (_zz_2250[31:0]        ), //i
    .dout    (fixTo_457_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_458 (
    .din     (_zz_2251[31:0]        ), //i
    .dout    (fixTo_458_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_459 (
    .din     (_zz_2252[31:0]        ), //i
    .dout    (fixTo_459_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_460 (
    .din     (_zz_2253[31:0]        ), //i
    .dout    (fixTo_460_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_461 (
    .din     (_zz_2254[31:0]        ), //i
    .dout    (fixTo_461_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_462 (
    .din     (_zz_2255[31:0]        ), //i
    .dout    (fixTo_462_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_463 (
    .din     (_zz_2256[31:0]        ), //i
    .dout    (fixTo_463_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_464 (
    .din     (_zz_2257[31:0]        ), //i
    .dout    (fixTo_464_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_465 (
    .din     (_zz_2258[31:0]        ), //i
    .dout    (fixTo_465_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_466 (
    .din     (_zz_2259[31:0]        ), //i
    .dout    (fixTo_466_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_467 (
    .din     (_zz_2260[31:0]        ), //i
    .dout    (fixTo_467_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_468 (
    .din     (_zz_2261[31:0]        ), //i
    .dout    (fixTo_468_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_469 (
    .din     (_zz_2262[31:0]        ), //i
    .dout    (fixTo_469_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_470 (
    .din     (_zz_2263[31:0]        ), //i
    .dout    (fixTo_470_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_471 (
    .din     (_zz_2264[31:0]        ), //i
    .dout    (fixTo_471_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_472 (
    .din     (_zz_2265[31:0]        ), //i
    .dout    (fixTo_472_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_473 (
    .din     (_zz_2266[31:0]        ), //i
    .dout    (fixTo_473_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_474 (
    .din     (_zz_2267[31:0]        ), //i
    .dout    (fixTo_474_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_475 (
    .din     (_zz_2268[31:0]        ), //i
    .dout    (fixTo_475_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_476 (
    .din     (_zz_2269[31:0]        ), //i
    .dout    (fixTo_476_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_477 (
    .din     (_zz_2270[31:0]        ), //i
    .dout    (fixTo_477_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_478 (
    .din     (_zz_2271[31:0]        ), //i
    .dout    (fixTo_478_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_479 (
    .din     (_zz_2272[31:0]        ), //i
    .dout    (fixTo_479_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_480 (
    .din     (_zz_2273[31:0]        ), //i
    .dout    (fixTo_480_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_481 (
    .din     (_zz_2274[31:0]        ), //i
    .dout    (fixTo_481_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_482 (
    .din     (_zz_2275[31:0]        ), //i
    .dout    (fixTo_482_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_483 (
    .din     (_zz_2276[31:0]        ), //i
    .dout    (fixTo_483_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_484 (
    .din     (_zz_2277[31:0]        ), //i
    .dout    (fixTo_484_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_485 (
    .din     (_zz_2278[31:0]        ), //i
    .dout    (fixTo_485_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_486 (
    .din     (_zz_2279[31:0]        ), //i
    .dout    (fixTo_486_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_487 (
    .din     (_zz_2280[31:0]        ), //i
    .dout    (fixTo_487_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_488 (
    .din     (_zz_2281[31:0]        ), //i
    .dout    (fixTo_488_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_489 (
    .din     (_zz_2282[31:0]        ), //i
    .dout    (fixTo_489_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_490 (
    .din     (_zz_2283[31:0]        ), //i
    .dout    (fixTo_490_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_491 (
    .din     (_zz_2284[31:0]        ), //i
    .dout    (fixTo_491_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_492 (
    .din     (_zz_2285[31:0]        ), //i
    .dout    (fixTo_492_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_493 (
    .din     (_zz_2286[31:0]        ), //i
    .dout    (fixTo_493_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_494 (
    .din     (_zz_2287[31:0]        ), //i
    .dout    (fixTo_494_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_495 (
    .din     (_zz_2288[31:0]        ), //i
    .dout    (fixTo_495_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_496 (
    .din     (_zz_2289[31:0]        ), //i
    .dout    (fixTo_496_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_497 (
    .din     (_zz_2290[31:0]        ), //i
    .dout    (fixTo_497_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_498 (
    .din     (_zz_2291[31:0]        ), //i
    .dout    (fixTo_498_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_499 (
    .din     (_zz_2292[31:0]        ), //i
    .dout    (fixTo_499_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_500 (
    .din     (_zz_2293[31:0]        ), //i
    .dout    (fixTo_500_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_501 (
    .din     (_zz_2294[31:0]        ), //i
    .dout    (fixTo_501_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_502 (
    .din     (_zz_2295[31:0]        ), //i
    .dout    (fixTo_502_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_503 (
    .din     (_zz_2296[31:0]        ), //i
    .dout    (fixTo_503_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_504 (
    .din     (_zz_2297[31:0]        ), //i
    .dout    (fixTo_504_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_505 (
    .din     (_zz_2298[31:0]        ), //i
    .dout    (fixTo_505_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_506 (
    .din     (_zz_2299[31:0]        ), //i
    .dout    (fixTo_506_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_507 (
    .din     (_zz_2300[31:0]        ), //i
    .dout    (fixTo_507_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_508 (
    .din     (_zz_2301[31:0]        ), //i
    .dout    (fixTo_508_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_509 (
    .din     (_zz_2302[31:0]        ), //i
    .dout    (fixTo_509_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_510 (
    .din     (_zz_2303[31:0]        ), //i
    .dout    (fixTo_510_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_511 (
    .din     (_zz_2304[31:0]        ), //i
    .dout    (fixTo_511_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_512 (
    .din     (_zz_2305[31:0]        ), //i
    .dout    (fixTo_512_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_513 (
    .din     (_zz_2306[31:0]        ), //i
    .dout    (fixTo_513_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_514 (
    .din     (_zz_2307[31:0]        ), //i
    .dout    (fixTo_514_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_515 (
    .din     (_zz_2308[31:0]        ), //i
    .dout    (fixTo_515_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_516 (
    .din     (_zz_2309[31:0]        ), //i
    .dout    (fixTo_516_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_517 (
    .din     (_zz_2310[31:0]        ), //i
    .dout    (fixTo_517_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_518 (
    .din     (_zz_2311[31:0]        ), //i
    .dout    (fixTo_518_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_519 (
    .din     (_zz_2312[31:0]        ), //i
    .dout    (fixTo_519_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_520 (
    .din     (_zz_2313[31:0]        ), //i
    .dout    (fixTo_520_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_521 (
    .din     (_zz_2314[31:0]        ), //i
    .dout    (fixTo_521_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_522 (
    .din     (_zz_2315[31:0]        ), //i
    .dout    (fixTo_522_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_523 (
    .din     (_zz_2316[31:0]        ), //i
    .dout    (fixTo_523_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_524 (
    .din     (_zz_2317[31:0]        ), //i
    .dout    (fixTo_524_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_525 (
    .din     (_zz_2318[31:0]        ), //i
    .dout    (fixTo_525_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_526 (
    .din     (_zz_2319[31:0]        ), //i
    .dout    (fixTo_526_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_527 (
    .din     (_zz_2320[31:0]        ), //i
    .dout    (fixTo_527_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_528 (
    .din     (_zz_2321[31:0]        ), //i
    .dout    (fixTo_528_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_529 (
    .din     (_zz_2322[31:0]        ), //i
    .dout    (fixTo_529_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_530 (
    .din     (_zz_2323[31:0]        ), //i
    .dout    (fixTo_530_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_531 (
    .din     (_zz_2324[31:0]        ), //i
    .dout    (fixTo_531_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_532 (
    .din     (_zz_2325[31:0]        ), //i
    .dout    (fixTo_532_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_533 (
    .din     (_zz_2326[31:0]        ), //i
    .dout    (fixTo_533_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_534 (
    .din     (_zz_2327[31:0]        ), //i
    .dout    (fixTo_534_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_535 (
    .din     (_zz_2328[31:0]        ), //i
    .dout    (fixTo_535_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_536 (
    .din     (_zz_2329[31:0]        ), //i
    .dout    (fixTo_536_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_537 (
    .din     (_zz_2330[31:0]        ), //i
    .dout    (fixTo_537_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_538 (
    .din     (_zz_2331[31:0]        ), //i
    .dout    (fixTo_538_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_539 (
    .din     (_zz_2332[31:0]        ), //i
    .dout    (fixTo_539_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_540 (
    .din     (_zz_2333[31:0]        ), //i
    .dout    (fixTo_540_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_541 (
    .din     (_zz_2334[31:0]        ), //i
    .dout    (fixTo_541_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_542 (
    .din     (_zz_2335[31:0]        ), //i
    .dout    (fixTo_542_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_543 (
    .din     (_zz_2336[31:0]        ), //i
    .dout    (fixTo_543_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_544 (
    .din     (_zz_2337[31:0]        ), //i
    .dout    (fixTo_544_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_545 (
    .din     (_zz_2338[31:0]        ), //i
    .dout    (fixTo_545_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_546 (
    .din     (_zz_2339[31:0]        ), //i
    .dout    (fixTo_546_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_547 (
    .din     (_zz_2340[31:0]        ), //i
    .dout    (fixTo_547_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_548 (
    .din     (_zz_2341[31:0]        ), //i
    .dout    (fixTo_548_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_549 (
    .din     (_zz_2342[31:0]        ), //i
    .dout    (fixTo_549_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_550 (
    .din     (_zz_2343[31:0]        ), //i
    .dout    (fixTo_550_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_551 (
    .din     (_zz_2344[31:0]        ), //i
    .dout    (fixTo_551_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_552 (
    .din     (_zz_2345[31:0]        ), //i
    .dout    (fixTo_552_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_553 (
    .din     (_zz_2346[31:0]        ), //i
    .dout    (fixTo_553_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_554 (
    .din     (_zz_2347[31:0]        ), //i
    .dout    (fixTo_554_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_555 (
    .din     (_zz_2348[31:0]        ), //i
    .dout    (fixTo_555_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_556 (
    .din     (_zz_2349[31:0]        ), //i
    .dout    (fixTo_556_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_557 (
    .din     (_zz_2350[31:0]        ), //i
    .dout    (fixTo_557_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_558 (
    .din     (_zz_2351[31:0]        ), //i
    .dout    (fixTo_558_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_559 (
    .din     (_zz_2352[31:0]        ), //i
    .dout    (fixTo_559_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_560 (
    .din     (_zz_2353[31:0]        ), //i
    .dout    (fixTo_560_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_561 (
    .din     (_zz_2354[31:0]        ), //i
    .dout    (fixTo_561_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_562 (
    .din     (_zz_2355[31:0]        ), //i
    .dout    (fixTo_562_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_563 (
    .din     (_zz_2356[31:0]        ), //i
    .dout    (fixTo_563_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_564 (
    .din     (_zz_2357[31:0]        ), //i
    .dout    (fixTo_564_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_565 (
    .din     (_zz_2358[31:0]        ), //i
    .dout    (fixTo_565_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_566 (
    .din     (_zz_2359[31:0]        ), //i
    .dout    (fixTo_566_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_567 (
    .din     (_zz_2360[31:0]        ), //i
    .dout    (fixTo_567_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_568 (
    .din     (_zz_2361[31:0]        ), //i
    .dout    (fixTo_568_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_569 (
    .din     (_zz_2362[31:0]        ), //i
    .dout    (fixTo_569_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_570 (
    .din     (_zz_2363[31:0]        ), //i
    .dout    (fixTo_570_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_571 (
    .din     (_zz_2364[31:0]        ), //i
    .dout    (fixTo_571_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_572 (
    .din     (_zz_2365[31:0]        ), //i
    .dout    (fixTo_572_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_573 (
    .din     (_zz_2366[31:0]        ), //i
    .dout    (fixTo_573_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_574 (
    .din     (_zz_2367[31:0]        ), //i
    .dout    (fixTo_574_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_575 (
    .din     (_zz_2368[31:0]        ), //i
    .dout    (fixTo_575_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_576 (
    .din     (_zz_2369[31:0]        ), //i
    .dout    (fixTo_576_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_577 (
    .din     (_zz_2370[31:0]        ), //i
    .dout    (fixTo_577_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_578 (
    .din     (_zz_2371[31:0]        ), //i
    .dout    (fixTo_578_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_579 (
    .din     (_zz_2372[31:0]        ), //i
    .dout    (fixTo_579_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_580 (
    .din     (_zz_2373[31:0]        ), //i
    .dout    (fixTo_580_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_581 (
    .din     (_zz_2374[31:0]        ), //i
    .dout    (fixTo_581_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_582 (
    .din     (_zz_2375[31:0]        ), //i
    .dout    (fixTo_582_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_583 (
    .din     (_zz_2376[31:0]        ), //i
    .dout    (fixTo_583_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_584 (
    .din     (_zz_2377[31:0]        ), //i
    .dout    (fixTo_584_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_585 (
    .din     (_zz_2378[31:0]        ), //i
    .dout    (fixTo_585_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_586 (
    .din     (_zz_2379[31:0]        ), //i
    .dout    (fixTo_586_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_587 (
    .din     (_zz_2380[31:0]        ), //i
    .dout    (fixTo_587_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_588 (
    .din     (_zz_2381[31:0]        ), //i
    .dout    (fixTo_588_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_589 (
    .din     (_zz_2382[31:0]        ), //i
    .dout    (fixTo_589_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_590 (
    .din     (_zz_2383[31:0]        ), //i
    .dout    (fixTo_590_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_591 (
    .din     (_zz_2384[31:0]        ), //i
    .dout    (fixTo_591_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_592 (
    .din     (_zz_2385[31:0]        ), //i
    .dout    (fixTo_592_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_593 (
    .din     (_zz_2386[31:0]        ), //i
    .dout    (fixTo_593_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_594 (
    .din     (_zz_2387[31:0]        ), //i
    .dout    (fixTo_594_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_595 (
    .din     (_zz_2388[31:0]        ), //i
    .dout    (fixTo_595_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_596 (
    .din     (_zz_2389[31:0]        ), //i
    .dout    (fixTo_596_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_597 (
    .din     (_zz_2390[31:0]        ), //i
    .dout    (fixTo_597_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_598 (
    .din     (_zz_2391[31:0]        ), //i
    .dout    (fixTo_598_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_599 (
    .din     (_zz_2392[31:0]        ), //i
    .dout    (fixTo_599_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_600 (
    .din     (_zz_2393[31:0]        ), //i
    .dout    (fixTo_600_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_601 (
    .din     (_zz_2394[31:0]        ), //i
    .dout    (fixTo_601_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_602 (
    .din     (_zz_2395[31:0]        ), //i
    .dout    (fixTo_602_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_603 (
    .din     (_zz_2396[31:0]        ), //i
    .dout    (fixTo_603_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_604 (
    .din     (_zz_2397[31:0]        ), //i
    .dout    (fixTo_604_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_605 (
    .din     (_zz_2398[31:0]        ), //i
    .dout    (fixTo_605_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_606 (
    .din     (_zz_2399[31:0]        ), //i
    .dout    (fixTo_606_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_607 (
    .din     (_zz_2400[31:0]        ), //i
    .dout    (fixTo_607_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_608 (
    .din     (_zz_2401[31:0]        ), //i
    .dout    (fixTo_608_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_609 (
    .din     (_zz_2402[31:0]        ), //i
    .dout    (fixTo_609_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_610 (
    .din     (_zz_2403[31:0]        ), //i
    .dout    (fixTo_610_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_611 (
    .din     (_zz_2404[31:0]        ), //i
    .dout    (fixTo_611_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_612 (
    .din     (_zz_2405[31:0]        ), //i
    .dout    (fixTo_612_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_613 (
    .din     (_zz_2406[31:0]        ), //i
    .dout    (fixTo_613_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_614 (
    .din     (_zz_2407[31:0]        ), //i
    .dout    (fixTo_614_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_615 (
    .din     (_zz_2408[31:0]        ), //i
    .dout    (fixTo_615_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_616 (
    .din     (_zz_2409[31:0]        ), //i
    .dout    (fixTo_616_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_617 (
    .din     (_zz_2410[31:0]        ), //i
    .dout    (fixTo_617_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_618 (
    .din     (_zz_2411[31:0]        ), //i
    .dout    (fixTo_618_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_619 (
    .din     (_zz_2412[31:0]        ), //i
    .dout    (fixTo_619_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_620 (
    .din     (_zz_2413[31:0]        ), //i
    .dout    (fixTo_620_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_621 (
    .din     (_zz_2414[31:0]        ), //i
    .dout    (fixTo_621_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_622 (
    .din     (_zz_2415[31:0]        ), //i
    .dout    (fixTo_622_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_623 (
    .din     (_zz_2416[31:0]        ), //i
    .dout    (fixTo_623_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_624 (
    .din     (_zz_2417[31:0]        ), //i
    .dout    (fixTo_624_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_625 (
    .din     (_zz_2418[31:0]        ), //i
    .dout    (fixTo_625_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_626 (
    .din     (_zz_2419[31:0]        ), //i
    .dout    (fixTo_626_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_627 (
    .din     (_zz_2420[31:0]        ), //i
    .dout    (fixTo_627_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_628 (
    .din     (_zz_2421[31:0]        ), //i
    .dout    (fixTo_628_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_629 (
    .din     (_zz_2422[31:0]        ), //i
    .dout    (fixTo_629_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_630 (
    .din     (_zz_2423[31:0]        ), //i
    .dout    (fixTo_630_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_631 (
    .din     (_zz_2424[31:0]        ), //i
    .dout    (fixTo_631_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_632 (
    .din     (_zz_2425[31:0]        ), //i
    .dout    (fixTo_632_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_633 (
    .din     (_zz_2426[31:0]        ), //i
    .dout    (fixTo_633_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_634 (
    .din     (_zz_2427[31:0]        ), //i
    .dout    (fixTo_634_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_635 (
    .din     (_zz_2428[31:0]        ), //i
    .dout    (fixTo_635_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_636 (
    .din     (_zz_2429[31:0]        ), //i
    .dout    (fixTo_636_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_637 (
    .din     (_zz_2430[31:0]        ), //i
    .dout    (fixTo_637_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_638 (
    .din     (_zz_2431[31:0]        ), //i
    .dout    (fixTo_638_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_639 (
    .din     (_zz_2432[31:0]        ), //i
    .dout    (fixTo_639_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_640 (
    .din     (_zz_2433[31:0]        ), //i
    .dout    (fixTo_640_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_641 (
    .din     (_zz_2434[31:0]        ), //i
    .dout    (fixTo_641_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_642 (
    .din     (_zz_2435[31:0]        ), //i
    .dout    (fixTo_642_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_643 (
    .din     (_zz_2436[31:0]        ), //i
    .dout    (fixTo_643_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_644 (
    .din     (_zz_2437[31:0]        ), //i
    .dout    (fixTo_644_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_645 (
    .din     (_zz_2438[31:0]        ), //i
    .dout    (fixTo_645_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_646 (
    .din     (_zz_2439[31:0]        ), //i
    .dout    (fixTo_646_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_647 (
    .din     (_zz_2440[31:0]        ), //i
    .dout    (fixTo_647_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_648 (
    .din     (_zz_2441[31:0]        ), //i
    .dout    (fixTo_648_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_649 (
    .din     (_zz_2442[31:0]        ), //i
    .dout    (fixTo_649_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_650 (
    .din     (_zz_2443[31:0]        ), //i
    .dout    (fixTo_650_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_651 (
    .din     (_zz_2444[31:0]        ), //i
    .dout    (fixTo_651_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_652 (
    .din     (_zz_2445[31:0]        ), //i
    .dout    (fixTo_652_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_653 (
    .din     (_zz_2446[31:0]        ), //i
    .dout    (fixTo_653_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_654 (
    .din     (_zz_2447[31:0]        ), //i
    .dout    (fixTo_654_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_655 (
    .din     (_zz_2448[31:0]        ), //i
    .dout    (fixTo_655_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_656 (
    .din     (_zz_2449[31:0]        ), //i
    .dout    (fixTo_656_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_657 (
    .din     (_zz_2450[31:0]        ), //i
    .dout    (fixTo_657_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_658 (
    .din     (_zz_2451[31:0]        ), //i
    .dout    (fixTo_658_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_659 (
    .din     (_zz_2452[31:0]        ), //i
    .dout    (fixTo_659_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_660 (
    .din     (_zz_2453[31:0]        ), //i
    .dout    (fixTo_660_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_661 (
    .din     (_zz_2454[31:0]        ), //i
    .dout    (fixTo_661_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_662 (
    .din     (_zz_2455[31:0]        ), //i
    .dout    (fixTo_662_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_663 (
    .din     (_zz_2456[31:0]        ), //i
    .dout    (fixTo_663_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_664 (
    .din     (_zz_2457[31:0]        ), //i
    .dout    (fixTo_664_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_665 (
    .din     (_zz_2458[31:0]        ), //i
    .dout    (fixTo_665_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_666 (
    .din     (_zz_2459[31:0]        ), //i
    .dout    (fixTo_666_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_667 (
    .din     (_zz_2460[31:0]        ), //i
    .dout    (fixTo_667_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_668 (
    .din     (_zz_2461[31:0]        ), //i
    .dout    (fixTo_668_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_669 (
    .din     (_zz_2462[31:0]        ), //i
    .dout    (fixTo_669_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_670 (
    .din     (_zz_2463[31:0]        ), //i
    .dout    (fixTo_670_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_671 (
    .din     (_zz_2464[31:0]        ), //i
    .dout    (fixTo_671_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_672 (
    .din     (_zz_2465[31:0]        ), //i
    .dout    (fixTo_672_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_673 (
    .din     (_zz_2466[31:0]        ), //i
    .dout    (fixTo_673_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_674 (
    .din     (_zz_2467[31:0]        ), //i
    .dout    (fixTo_674_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_675 (
    .din     (_zz_2468[31:0]        ), //i
    .dout    (fixTo_675_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_676 (
    .din     (_zz_2469[31:0]        ), //i
    .dout    (fixTo_676_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_677 (
    .din     (_zz_2470[31:0]        ), //i
    .dout    (fixTo_677_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_678 (
    .din     (_zz_2471[31:0]        ), //i
    .dout    (fixTo_678_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_679 (
    .din     (_zz_2472[31:0]        ), //i
    .dout    (fixTo_679_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_680 (
    .din     (_zz_2473[31:0]        ), //i
    .dout    (fixTo_680_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_681 (
    .din     (_zz_2474[31:0]        ), //i
    .dout    (fixTo_681_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_682 (
    .din     (_zz_2475[31:0]        ), //i
    .dout    (fixTo_682_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_683 (
    .din     (_zz_2476[31:0]        ), //i
    .dout    (fixTo_683_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_684 (
    .din     (_zz_2477[31:0]        ), //i
    .dout    (fixTo_684_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_685 (
    .din     (_zz_2478[31:0]        ), //i
    .dout    (fixTo_685_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_686 (
    .din     (_zz_2479[31:0]        ), //i
    .dout    (fixTo_686_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_687 (
    .din     (_zz_2480[31:0]        ), //i
    .dout    (fixTo_687_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_688 (
    .din     (_zz_2481[31:0]        ), //i
    .dout    (fixTo_688_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_689 (
    .din     (_zz_2482[31:0]        ), //i
    .dout    (fixTo_689_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_690 (
    .din     (_zz_2483[31:0]        ), //i
    .dout    (fixTo_690_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_691 (
    .din     (_zz_2484[31:0]        ), //i
    .dout    (fixTo_691_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_692 (
    .din     (_zz_2485[31:0]        ), //i
    .dout    (fixTo_692_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_693 (
    .din     (_zz_2486[31:0]        ), //i
    .dout    (fixTo_693_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_694 (
    .din     (_zz_2487[31:0]        ), //i
    .dout    (fixTo_694_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_695 (
    .din     (_zz_2488[31:0]        ), //i
    .dout    (fixTo_695_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_696 (
    .din     (_zz_2489[31:0]        ), //i
    .dout    (fixTo_696_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_697 (
    .din     (_zz_2490[31:0]        ), //i
    .dout    (fixTo_697_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_698 (
    .din     (_zz_2491[31:0]        ), //i
    .dout    (fixTo_698_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_699 (
    .din     (_zz_2492[31:0]        ), //i
    .dout    (fixTo_699_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_700 (
    .din     (_zz_2493[31:0]        ), //i
    .dout    (fixTo_700_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_701 (
    .din     (_zz_2494[31:0]        ), //i
    .dout    (fixTo_701_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_702 (
    .din     (_zz_2495[31:0]        ), //i
    .dout    (fixTo_702_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_703 (
    .din     (_zz_2496[31:0]        ), //i
    .dout    (fixTo_703_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_704 (
    .din     (_zz_2497[31:0]        ), //i
    .dout    (fixTo_704_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_705 (
    .din     (_zz_2498[31:0]        ), //i
    .dout    (fixTo_705_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_706 (
    .din     (_zz_2499[31:0]        ), //i
    .dout    (fixTo_706_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_707 (
    .din     (_zz_2500[31:0]        ), //i
    .dout    (fixTo_707_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_708 (
    .din     (_zz_2501[31:0]        ), //i
    .dout    (fixTo_708_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_709 (
    .din     (_zz_2502[31:0]        ), //i
    .dout    (fixTo_709_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_710 (
    .din     (_zz_2503[31:0]        ), //i
    .dout    (fixTo_710_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_711 (
    .din     (_zz_2504[31:0]        ), //i
    .dout    (fixTo_711_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_712 (
    .din     (_zz_2505[31:0]        ), //i
    .dout    (fixTo_712_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_713 (
    .din     (_zz_2506[31:0]        ), //i
    .dout    (fixTo_713_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_714 (
    .din     (_zz_2507[31:0]        ), //i
    .dout    (fixTo_714_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_715 (
    .din     (_zz_2508[31:0]        ), //i
    .dout    (fixTo_715_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_716 (
    .din     (_zz_2509[31:0]        ), //i
    .dout    (fixTo_716_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_717 (
    .din     (_zz_2510[31:0]        ), //i
    .dout    (fixTo_717_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_718 (
    .din     (_zz_2511[31:0]        ), //i
    .dout    (fixTo_718_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_719 (
    .din     (_zz_2512[31:0]        ), //i
    .dout    (fixTo_719_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_720 (
    .din     (_zz_2513[31:0]        ), //i
    .dout    (fixTo_720_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_721 (
    .din     (_zz_2514[31:0]        ), //i
    .dout    (fixTo_721_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_722 (
    .din     (_zz_2515[31:0]        ), //i
    .dout    (fixTo_722_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_723 (
    .din     (_zz_2516[31:0]        ), //i
    .dout    (fixTo_723_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_724 (
    .din     (_zz_2517[31:0]        ), //i
    .dout    (fixTo_724_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_725 (
    .din     (_zz_2518[31:0]        ), //i
    .dout    (fixTo_725_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_726 (
    .din     (_zz_2519[31:0]        ), //i
    .dout    (fixTo_726_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_727 (
    .din     (_zz_2520[31:0]        ), //i
    .dout    (fixTo_727_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_728 (
    .din     (_zz_2521[31:0]        ), //i
    .dout    (fixTo_728_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_729 (
    .din     (_zz_2522[31:0]        ), //i
    .dout    (fixTo_729_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_730 (
    .din     (_zz_2523[31:0]        ), //i
    .dout    (fixTo_730_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_731 (
    .din     (_zz_2524[31:0]        ), //i
    .dout    (fixTo_731_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_732 (
    .din     (_zz_2525[31:0]        ), //i
    .dout    (fixTo_732_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_733 (
    .din     (_zz_2526[31:0]        ), //i
    .dout    (fixTo_733_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_734 (
    .din     (_zz_2527[31:0]        ), //i
    .dout    (fixTo_734_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_735 (
    .din     (_zz_2528[31:0]        ), //i
    .dout    (fixTo_735_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_736 (
    .din     (_zz_2529[31:0]        ), //i
    .dout    (fixTo_736_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_737 (
    .din     (_zz_2530[31:0]        ), //i
    .dout    (fixTo_737_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_738 (
    .din     (_zz_2531[31:0]        ), //i
    .dout    (fixTo_738_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_739 (
    .din     (_zz_2532[31:0]        ), //i
    .dout    (fixTo_739_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_740 (
    .din     (_zz_2533[31:0]        ), //i
    .dout    (fixTo_740_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_741 (
    .din     (_zz_2534[31:0]        ), //i
    .dout    (fixTo_741_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_742 (
    .din     (_zz_2535[31:0]        ), //i
    .dout    (fixTo_742_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_743 (
    .din     (_zz_2536[31:0]        ), //i
    .dout    (fixTo_743_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_744 (
    .din     (_zz_2537[31:0]        ), //i
    .dout    (fixTo_744_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_745 (
    .din     (_zz_2538[31:0]        ), //i
    .dout    (fixTo_745_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_746 (
    .din     (_zz_2539[31:0]        ), //i
    .dout    (fixTo_746_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_747 (
    .din     (_zz_2540[31:0]        ), //i
    .dout    (fixTo_747_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_748 (
    .din     (_zz_2541[31:0]        ), //i
    .dout    (fixTo_748_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_749 (
    .din     (_zz_2542[31:0]        ), //i
    .dout    (fixTo_749_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_750 (
    .din     (_zz_2543[31:0]        ), //i
    .dout    (fixTo_750_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_751 (
    .din     (_zz_2544[31:0]        ), //i
    .dout    (fixTo_751_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_752 (
    .din     (_zz_2545[31:0]        ), //i
    .dout    (fixTo_752_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_753 (
    .din     (_zz_2546[31:0]        ), //i
    .dout    (fixTo_753_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_754 (
    .din     (_zz_2547[31:0]        ), //i
    .dout    (fixTo_754_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_755 (
    .din     (_zz_2548[31:0]        ), //i
    .dout    (fixTo_755_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_756 (
    .din     (_zz_2549[31:0]        ), //i
    .dout    (fixTo_756_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_757 (
    .din     (_zz_2550[31:0]        ), //i
    .dout    (fixTo_757_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_758 (
    .din     (_zz_2551[31:0]        ), //i
    .dout    (fixTo_758_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_759 (
    .din     (_zz_2552[31:0]        ), //i
    .dout    (fixTo_759_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_760 (
    .din     (_zz_2553[31:0]        ), //i
    .dout    (fixTo_760_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_761 (
    .din     (_zz_2554[31:0]        ), //i
    .dout    (fixTo_761_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_762 (
    .din     (_zz_2555[31:0]        ), //i
    .dout    (fixTo_762_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_763 (
    .din     (_zz_2556[31:0]        ), //i
    .dout    (fixTo_763_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_764 (
    .din     (_zz_2557[31:0]        ), //i
    .dout    (fixTo_764_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_765 (
    .din     (_zz_2558[31:0]        ), //i
    .dout    (fixTo_765_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_766 (
    .din     (_zz_2559[31:0]        ), //i
    .dout    (fixTo_766_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_767 (
    .din     (_zz_2560[31:0]        ), //i
    .dout    (fixTo_767_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_768 (
    .din     (_zz_2561[31:0]        ), //i
    .dout    (fixTo_768_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_769 (
    .din     (_zz_2562[31:0]        ), //i
    .dout    (fixTo_769_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_770 (
    .din     (_zz_2563[31:0]        ), //i
    .dout    (fixTo_770_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_771 (
    .din     (_zz_2564[31:0]        ), //i
    .dout    (fixTo_771_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_772 (
    .din     (_zz_2565[31:0]        ), //i
    .dout    (fixTo_772_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_773 (
    .din     (_zz_2566[31:0]        ), //i
    .dout    (fixTo_773_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_774 (
    .din     (_zz_2567[31:0]        ), //i
    .dout    (fixTo_774_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_775 (
    .din     (_zz_2568[31:0]        ), //i
    .dout    (fixTo_775_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_776 (
    .din     (_zz_2569[31:0]        ), //i
    .dout    (fixTo_776_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_777 (
    .din     (_zz_2570[31:0]        ), //i
    .dout    (fixTo_777_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_778 (
    .din     (_zz_2571[31:0]        ), //i
    .dout    (fixTo_778_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_779 (
    .din     (_zz_2572[31:0]        ), //i
    .dout    (fixTo_779_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_780 (
    .din     (_zz_2573[31:0]        ), //i
    .dout    (fixTo_780_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_781 (
    .din     (_zz_2574[31:0]        ), //i
    .dout    (fixTo_781_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_782 (
    .din     (_zz_2575[31:0]        ), //i
    .dout    (fixTo_782_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_783 (
    .din     (_zz_2576[31:0]        ), //i
    .dout    (fixTo_783_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_784 (
    .din     (_zz_2577[31:0]        ), //i
    .dout    (fixTo_784_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_785 (
    .din     (_zz_2578[31:0]        ), //i
    .dout    (fixTo_785_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_786 (
    .din     (_zz_2579[31:0]        ), //i
    .dout    (fixTo_786_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_787 (
    .din     (_zz_2580[31:0]        ), //i
    .dout    (fixTo_787_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_788 (
    .din     (_zz_2581[31:0]        ), //i
    .dout    (fixTo_788_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_789 (
    .din     (_zz_2582[31:0]        ), //i
    .dout    (fixTo_789_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_790 (
    .din     (_zz_2583[31:0]        ), //i
    .dout    (fixTo_790_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_791 (
    .din     (_zz_2584[31:0]        ), //i
    .dout    (fixTo_791_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_792 (
    .din     (_zz_2585[31:0]        ), //i
    .dout    (fixTo_792_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_793 (
    .din     (_zz_2586[31:0]        ), //i
    .dout    (fixTo_793_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_794 (
    .din     (_zz_2587[31:0]        ), //i
    .dout    (fixTo_794_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_795 (
    .din     (_zz_2588[31:0]        ), //i
    .dout    (fixTo_795_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_796 (
    .din     (_zz_2589[31:0]        ), //i
    .dout    (fixTo_796_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_797 (
    .din     (_zz_2590[31:0]        ), //i
    .dout    (fixTo_797_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_798 (
    .din     (_zz_2591[31:0]        ), //i
    .dout    (fixTo_798_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_799 (
    .din     (_zz_2592[31:0]        ), //i
    .dout    (fixTo_799_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_800 (
    .din     (_zz_2593[31:0]        ), //i
    .dout    (fixTo_800_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_801 (
    .din     (_zz_2594[31:0]        ), //i
    .dout    (fixTo_801_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_802 (
    .din     (_zz_2595[31:0]        ), //i
    .dout    (fixTo_802_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_803 (
    .din     (_zz_2596[31:0]        ), //i
    .dout    (fixTo_803_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_804 (
    .din     (_zz_2597[31:0]        ), //i
    .dout    (fixTo_804_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_805 (
    .din     (_zz_2598[31:0]        ), //i
    .dout    (fixTo_805_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_806 (
    .din     (_zz_2599[31:0]        ), //i
    .dout    (fixTo_806_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_807 (
    .din     (_zz_2600[31:0]        ), //i
    .dout    (fixTo_807_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_808 (
    .din     (_zz_2601[31:0]        ), //i
    .dout    (fixTo_808_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_809 (
    .din     (_zz_2602[31:0]        ), //i
    .dout    (fixTo_809_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_810 (
    .din     (_zz_2603[31:0]        ), //i
    .dout    (fixTo_810_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_811 (
    .din     (_zz_2604[31:0]        ), //i
    .dout    (fixTo_811_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_812 (
    .din     (_zz_2605[31:0]        ), //i
    .dout    (fixTo_812_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_813 (
    .din     (_zz_2606[31:0]        ), //i
    .dout    (fixTo_813_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_814 (
    .din     (_zz_2607[31:0]        ), //i
    .dout    (fixTo_814_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_815 (
    .din     (_zz_2608[31:0]        ), //i
    .dout    (fixTo_815_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_816 (
    .din     (_zz_2609[31:0]        ), //i
    .dout    (fixTo_816_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_817 (
    .din     (_zz_2610[31:0]        ), //i
    .dout    (fixTo_817_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_818 (
    .din     (_zz_2611[31:0]        ), //i
    .dout    (fixTo_818_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_819 (
    .din     (_zz_2612[31:0]        ), //i
    .dout    (fixTo_819_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_820 (
    .din     (_zz_2613[31:0]        ), //i
    .dout    (fixTo_820_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_821 (
    .din     (_zz_2614[31:0]        ), //i
    .dout    (fixTo_821_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_822 (
    .din     (_zz_2615[31:0]        ), //i
    .dout    (fixTo_822_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_823 (
    .din     (_zz_2616[31:0]        ), //i
    .dout    (fixTo_823_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_824 (
    .din     (_zz_2617[31:0]        ), //i
    .dout    (fixTo_824_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_825 (
    .din     (_zz_2618[31:0]        ), //i
    .dout    (fixTo_825_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_826 (
    .din     (_zz_2619[31:0]        ), //i
    .dout    (fixTo_826_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_827 (
    .din     (_zz_2620[31:0]        ), //i
    .dout    (fixTo_827_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_828 (
    .din     (_zz_2621[31:0]        ), //i
    .dout    (fixTo_828_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_829 (
    .din     (_zz_2622[31:0]        ), //i
    .dout    (fixTo_829_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_830 (
    .din     (_zz_2623[31:0]        ), //i
    .dout    (fixTo_830_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_831 (
    .din     (_zz_2624[31:0]        ), //i
    .dout    (fixTo_831_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_832 (
    .din     (_zz_2625[31:0]        ), //i
    .dout    (fixTo_832_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_833 (
    .din     (_zz_2626[31:0]        ), //i
    .dout    (fixTo_833_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_834 (
    .din     (_zz_2627[31:0]        ), //i
    .dout    (fixTo_834_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_835 (
    .din     (_zz_2628[31:0]        ), //i
    .dout    (fixTo_835_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_836 (
    .din     (_zz_2629[31:0]        ), //i
    .dout    (fixTo_836_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_837 (
    .din     (_zz_2630[31:0]        ), //i
    .dout    (fixTo_837_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_838 (
    .din     (_zz_2631[31:0]        ), //i
    .dout    (fixTo_838_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_839 (
    .din     (_zz_2632[31:0]        ), //i
    .dout    (fixTo_839_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_840 (
    .din     (_zz_2633[31:0]        ), //i
    .dout    (fixTo_840_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_841 (
    .din     (_zz_2634[31:0]        ), //i
    .dout    (fixTo_841_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_842 (
    .din     (_zz_2635[31:0]        ), //i
    .dout    (fixTo_842_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_843 (
    .din     (_zz_2636[31:0]        ), //i
    .dout    (fixTo_843_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_844 (
    .din     (_zz_2637[31:0]        ), //i
    .dout    (fixTo_844_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_845 (
    .din     (_zz_2638[31:0]        ), //i
    .dout    (fixTo_845_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_846 (
    .din     (_zz_2639[31:0]        ), //i
    .dout    (fixTo_846_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_847 (
    .din     (_zz_2640[31:0]        ), //i
    .dout    (fixTo_847_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_848 (
    .din     (_zz_2641[31:0]        ), //i
    .dout    (fixTo_848_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_849 (
    .din     (_zz_2642[31:0]        ), //i
    .dout    (fixTo_849_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_850 (
    .din     (_zz_2643[31:0]        ), //i
    .dout    (fixTo_850_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_851 (
    .din     (_zz_2644[31:0]        ), //i
    .dout    (fixTo_851_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_852 (
    .din     (_zz_2645[31:0]        ), //i
    .dout    (fixTo_852_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_853 (
    .din     (_zz_2646[31:0]        ), //i
    .dout    (fixTo_853_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_854 (
    .din     (_zz_2647[31:0]        ), //i
    .dout    (fixTo_854_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_855 (
    .din     (_zz_2648[31:0]        ), //i
    .dout    (fixTo_855_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_856 (
    .din     (_zz_2649[31:0]        ), //i
    .dout    (fixTo_856_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_857 (
    .din     (_zz_2650[31:0]        ), //i
    .dout    (fixTo_857_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_858 (
    .din     (_zz_2651[31:0]        ), //i
    .dout    (fixTo_858_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_859 (
    .din     (_zz_2652[31:0]        ), //i
    .dout    (fixTo_859_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_860 (
    .din     (_zz_2653[31:0]        ), //i
    .dout    (fixTo_860_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_861 (
    .din     (_zz_2654[31:0]        ), //i
    .dout    (fixTo_861_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_862 (
    .din     (_zz_2655[31:0]        ), //i
    .dout    (fixTo_862_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_863 (
    .din     (_zz_2656[31:0]        ), //i
    .dout    (fixTo_863_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_864 (
    .din     (_zz_2657[31:0]        ), //i
    .dout    (fixTo_864_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_865 (
    .din     (_zz_2658[31:0]        ), //i
    .dout    (fixTo_865_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_866 (
    .din     (_zz_2659[31:0]        ), //i
    .dout    (fixTo_866_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_867 (
    .din     (_zz_2660[31:0]        ), //i
    .dout    (fixTo_867_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_868 (
    .din     (_zz_2661[31:0]        ), //i
    .dout    (fixTo_868_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_869 (
    .din     (_zz_2662[31:0]        ), //i
    .dout    (fixTo_869_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_870 (
    .din     (_zz_2663[31:0]        ), //i
    .dout    (fixTo_870_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_871 (
    .din     (_zz_2664[31:0]        ), //i
    .dout    (fixTo_871_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_872 (
    .din     (_zz_2665[31:0]        ), //i
    .dout    (fixTo_872_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_873 (
    .din     (_zz_2666[31:0]        ), //i
    .dout    (fixTo_873_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_874 (
    .din     (_zz_2667[31:0]        ), //i
    .dout    (fixTo_874_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_875 (
    .din     (_zz_2668[31:0]        ), //i
    .dout    (fixTo_875_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_876 (
    .din     (_zz_2669[31:0]        ), //i
    .dout    (fixTo_876_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_877 (
    .din     (_zz_2670[31:0]        ), //i
    .dout    (fixTo_877_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_878 (
    .din     (_zz_2671[31:0]        ), //i
    .dout    (fixTo_878_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_879 (
    .din     (_zz_2672[31:0]        ), //i
    .dout    (fixTo_879_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_880 (
    .din     (_zz_2673[31:0]        ), //i
    .dout    (fixTo_880_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_881 (
    .din     (_zz_2674[31:0]        ), //i
    .dout    (fixTo_881_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_882 (
    .din     (_zz_2675[31:0]        ), //i
    .dout    (fixTo_882_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_883 (
    .din     (_zz_2676[31:0]        ), //i
    .dout    (fixTo_883_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_884 (
    .din     (_zz_2677[31:0]        ), //i
    .dout    (fixTo_884_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_885 (
    .din     (_zz_2678[31:0]        ), //i
    .dout    (fixTo_885_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_886 (
    .din     (_zz_2679[31:0]        ), //i
    .dout    (fixTo_886_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_887 (
    .din     (_zz_2680[31:0]        ), //i
    .dout    (fixTo_887_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_888 (
    .din     (_zz_2681[31:0]        ), //i
    .dout    (fixTo_888_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_889 (
    .din     (_zz_2682[31:0]        ), //i
    .dout    (fixTo_889_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_890 (
    .din     (_zz_2683[31:0]        ), //i
    .dout    (fixTo_890_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_891 (
    .din     (_zz_2684[31:0]        ), //i
    .dout    (fixTo_891_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_892 (
    .din     (_zz_2685[31:0]        ), //i
    .dout    (fixTo_892_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_893 (
    .din     (_zz_2686[31:0]        ), //i
    .dout    (fixTo_893_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_894 (
    .din     (_zz_2687[31:0]        ), //i
    .dout    (fixTo_894_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_895 (
    .din     (_zz_2688[31:0]        ), //i
    .dout    (fixTo_895_dout[15:0]  )  //o
  );
  assign twiddle_factor_table_0_real = 16'h0100;
  assign twiddle_factor_table_0_imag = 16'h0;
  assign twiddle_factor_table_1_real = 16'h0100;
  assign twiddle_factor_table_1_imag = 16'h0;
  assign twiddle_factor_table_2_real = 16'h0;
  assign twiddle_factor_table_2_imag = 16'hff00;
  assign twiddle_factor_table_3_real = 16'h0100;
  assign twiddle_factor_table_3_imag = 16'h0;
  assign twiddle_factor_table_4_real = 16'h00b5;
  assign twiddle_factor_table_4_imag = 16'hff4b;
  assign twiddle_factor_table_5_real = 16'h0;
  assign twiddle_factor_table_5_imag = 16'hff00;
  assign twiddle_factor_table_6_real = 16'hff4b;
  assign twiddle_factor_table_6_imag = 16'hff4b;
  assign twiddle_factor_table_7_real = 16'h0100;
  assign twiddle_factor_table_7_imag = 16'h0;
  assign twiddle_factor_table_8_real = 16'h00ec;
  assign twiddle_factor_table_8_imag = 16'hff9f;
  assign twiddle_factor_table_9_real = 16'h00b5;
  assign twiddle_factor_table_9_imag = 16'hff4b;
  assign twiddle_factor_table_10_real = 16'h0061;
  assign twiddle_factor_table_10_imag = 16'hff14;
  assign twiddle_factor_table_11_real = 16'h0;
  assign twiddle_factor_table_11_imag = 16'hff00;
  assign twiddle_factor_table_12_real = 16'hff9f;
  assign twiddle_factor_table_12_imag = 16'hff14;
  assign twiddle_factor_table_13_real = 16'hff4b;
  assign twiddle_factor_table_13_imag = 16'hff4b;
  assign twiddle_factor_table_14_real = 16'hff14;
  assign twiddle_factor_table_14_imag = 16'hff9f;
  assign twiddle_factor_table_15_real = 16'h0100;
  assign twiddle_factor_table_15_imag = 16'h0;
  assign twiddle_factor_table_16_real = 16'h00fb;
  assign twiddle_factor_table_16_imag = 16'hffcf;
  assign twiddle_factor_table_17_real = 16'h00ec;
  assign twiddle_factor_table_17_imag = 16'hff9f;
  assign twiddle_factor_table_18_real = 16'h00d4;
  assign twiddle_factor_table_18_imag = 16'hff72;
  assign twiddle_factor_table_19_real = 16'h00b5;
  assign twiddle_factor_table_19_imag = 16'hff4b;
  assign twiddle_factor_table_20_real = 16'h008e;
  assign twiddle_factor_table_20_imag = 16'hff2c;
  assign twiddle_factor_table_21_real = 16'h0061;
  assign twiddle_factor_table_21_imag = 16'hff14;
  assign twiddle_factor_table_22_real = 16'h0031;
  assign twiddle_factor_table_22_imag = 16'hff05;
  assign twiddle_factor_table_23_real = 16'h0;
  assign twiddle_factor_table_23_imag = 16'hff00;
  assign twiddle_factor_table_24_real = 16'hffcf;
  assign twiddle_factor_table_24_imag = 16'hff05;
  assign twiddle_factor_table_25_real = 16'hff9f;
  assign twiddle_factor_table_25_imag = 16'hff14;
  assign twiddle_factor_table_26_real = 16'hff72;
  assign twiddle_factor_table_26_imag = 16'hff2c;
  assign twiddle_factor_table_27_real = 16'hff4b;
  assign twiddle_factor_table_27_imag = 16'hff4b;
  assign twiddle_factor_table_28_real = 16'hff2c;
  assign twiddle_factor_table_28_imag = 16'hff72;
  assign twiddle_factor_table_29_real = 16'hff14;
  assign twiddle_factor_table_29_imag = 16'hff9f;
  assign twiddle_factor_table_30_real = 16'hff05;
  assign twiddle_factor_table_30_imag = 16'hffcf;
  assign twiddle_factor_table_31_real = 16'h0100;
  assign twiddle_factor_table_31_imag = 16'h0;
  assign twiddle_factor_table_32_real = 16'h00fe;
  assign twiddle_factor_table_32_imag = 16'hffe7;
  assign twiddle_factor_table_33_real = 16'h00fb;
  assign twiddle_factor_table_33_imag = 16'hffcf;
  assign twiddle_factor_table_34_real = 16'h00f4;
  assign twiddle_factor_table_34_imag = 16'hffb6;
  assign twiddle_factor_table_35_real = 16'h00ec;
  assign twiddle_factor_table_35_imag = 16'hff9f;
  assign twiddle_factor_table_36_real = 16'h00e1;
  assign twiddle_factor_table_36_imag = 16'hff88;
  assign twiddle_factor_table_37_real = 16'h00d4;
  assign twiddle_factor_table_37_imag = 16'hff72;
  assign twiddle_factor_table_38_real = 16'h00c5;
  assign twiddle_factor_table_38_imag = 16'hff5e;
  assign twiddle_factor_table_39_real = 16'h00b5;
  assign twiddle_factor_table_39_imag = 16'hff4b;
  assign twiddle_factor_table_40_real = 16'h00a2;
  assign twiddle_factor_table_40_imag = 16'hff3b;
  assign twiddle_factor_table_41_real = 16'h008e;
  assign twiddle_factor_table_41_imag = 16'hff2c;
  assign twiddle_factor_table_42_real = 16'h0078;
  assign twiddle_factor_table_42_imag = 16'hff1f;
  assign twiddle_factor_table_43_real = 16'h0061;
  assign twiddle_factor_table_43_imag = 16'hff14;
  assign twiddle_factor_table_44_real = 16'h004a;
  assign twiddle_factor_table_44_imag = 16'hff0c;
  assign twiddle_factor_table_45_real = 16'h0031;
  assign twiddle_factor_table_45_imag = 16'hff05;
  assign twiddle_factor_table_46_real = 16'h0019;
  assign twiddle_factor_table_46_imag = 16'hff02;
  assign twiddle_factor_table_47_real = 16'h0;
  assign twiddle_factor_table_47_imag = 16'hff00;
  assign twiddle_factor_table_48_real = 16'hffe7;
  assign twiddle_factor_table_48_imag = 16'hff02;
  assign twiddle_factor_table_49_real = 16'hffcf;
  assign twiddle_factor_table_49_imag = 16'hff05;
  assign twiddle_factor_table_50_real = 16'hffb6;
  assign twiddle_factor_table_50_imag = 16'hff0c;
  assign twiddle_factor_table_51_real = 16'hff9f;
  assign twiddle_factor_table_51_imag = 16'hff14;
  assign twiddle_factor_table_52_real = 16'hff88;
  assign twiddle_factor_table_52_imag = 16'hff1f;
  assign twiddle_factor_table_53_real = 16'hff72;
  assign twiddle_factor_table_53_imag = 16'hff2c;
  assign twiddle_factor_table_54_real = 16'hff5e;
  assign twiddle_factor_table_54_imag = 16'hff3b;
  assign twiddle_factor_table_55_real = 16'hff4b;
  assign twiddle_factor_table_55_imag = 16'hff4b;
  assign twiddle_factor_table_56_real = 16'hff3b;
  assign twiddle_factor_table_56_imag = 16'hff5e;
  assign twiddle_factor_table_57_real = 16'hff2c;
  assign twiddle_factor_table_57_imag = 16'hff72;
  assign twiddle_factor_table_58_real = 16'hff1f;
  assign twiddle_factor_table_58_imag = 16'hff88;
  assign twiddle_factor_table_59_real = 16'hff14;
  assign twiddle_factor_table_59_imag = 16'hff9f;
  assign twiddle_factor_table_60_real = 16'hff0c;
  assign twiddle_factor_table_60_imag = 16'hffb6;
  assign twiddle_factor_table_61_real = 16'hff05;
  assign twiddle_factor_table_61_imag = 16'hffcf;
  assign twiddle_factor_table_62_real = 16'hff02;
  assign twiddle_factor_table_62_imag = 16'hffe7;
  assign twiddle_factor_table_63_real = 16'h0100;
  assign twiddle_factor_table_63_imag = 16'h0;
  assign twiddle_factor_table_64_real = 16'h00ff;
  assign twiddle_factor_table_64_imag = 16'hfff4;
  assign twiddle_factor_table_65_real = 16'h00fe;
  assign twiddle_factor_table_65_imag = 16'hffe7;
  assign twiddle_factor_table_66_real = 16'h00fd;
  assign twiddle_factor_table_66_imag = 16'hffdb;
  assign twiddle_factor_table_67_real = 16'h00fb;
  assign twiddle_factor_table_67_imag = 16'hffcf;
  assign twiddle_factor_table_68_real = 16'h00f8;
  assign twiddle_factor_table_68_imag = 16'hffc2;
  assign twiddle_factor_table_69_real = 16'h00f4;
  assign twiddle_factor_table_69_imag = 16'hffb6;
  assign twiddle_factor_table_70_real = 16'h00f1;
  assign twiddle_factor_table_70_imag = 16'hffaa;
  assign twiddle_factor_table_71_real = 16'h00ec;
  assign twiddle_factor_table_71_imag = 16'hff9f;
  assign twiddle_factor_table_72_real = 16'h00e7;
  assign twiddle_factor_table_72_imag = 16'hff93;
  assign twiddle_factor_table_73_real = 16'h00e1;
  assign twiddle_factor_table_73_imag = 16'hff88;
  assign twiddle_factor_table_74_real = 16'h00db;
  assign twiddle_factor_table_74_imag = 16'hff7d;
  assign twiddle_factor_table_75_real = 16'h00d4;
  assign twiddle_factor_table_75_imag = 16'hff72;
  assign twiddle_factor_table_76_real = 16'h00cd;
  assign twiddle_factor_table_76_imag = 16'hff68;
  assign twiddle_factor_table_77_real = 16'h00c5;
  assign twiddle_factor_table_77_imag = 16'hff5e;
  assign twiddle_factor_table_78_real = 16'h00bd;
  assign twiddle_factor_table_78_imag = 16'hff55;
  assign twiddle_factor_table_79_real = 16'h00b5;
  assign twiddle_factor_table_79_imag = 16'hff4b;
  assign twiddle_factor_table_80_real = 16'h00ab;
  assign twiddle_factor_table_80_imag = 16'hff43;
  assign twiddle_factor_table_81_real = 16'h00a2;
  assign twiddle_factor_table_81_imag = 16'hff3b;
  assign twiddle_factor_table_82_real = 16'h0098;
  assign twiddle_factor_table_82_imag = 16'hff33;
  assign twiddle_factor_table_83_real = 16'h008e;
  assign twiddle_factor_table_83_imag = 16'hff2c;
  assign twiddle_factor_table_84_real = 16'h0083;
  assign twiddle_factor_table_84_imag = 16'hff25;
  assign twiddle_factor_table_85_real = 16'h0078;
  assign twiddle_factor_table_85_imag = 16'hff1f;
  assign twiddle_factor_table_86_real = 16'h006d;
  assign twiddle_factor_table_86_imag = 16'hff19;
  assign twiddle_factor_table_87_real = 16'h0061;
  assign twiddle_factor_table_87_imag = 16'hff14;
  assign twiddle_factor_table_88_real = 16'h0056;
  assign twiddle_factor_table_88_imag = 16'hff0f;
  assign twiddle_factor_table_89_real = 16'h004a;
  assign twiddle_factor_table_89_imag = 16'hff0c;
  assign twiddle_factor_table_90_real = 16'h003e;
  assign twiddle_factor_table_90_imag = 16'hff08;
  assign twiddle_factor_table_91_real = 16'h0031;
  assign twiddle_factor_table_91_imag = 16'hff05;
  assign twiddle_factor_table_92_real = 16'h0025;
  assign twiddle_factor_table_92_imag = 16'hff03;
  assign twiddle_factor_table_93_real = 16'h0019;
  assign twiddle_factor_table_93_imag = 16'hff02;
  assign twiddle_factor_table_94_real = 16'h000c;
  assign twiddle_factor_table_94_imag = 16'hff01;
  assign twiddle_factor_table_95_real = 16'h0;
  assign twiddle_factor_table_95_imag = 16'hff00;
  assign twiddle_factor_table_96_real = 16'hfff4;
  assign twiddle_factor_table_96_imag = 16'hff01;
  assign twiddle_factor_table_97_real = 16'hffe7;
  assign twiddle_factor_table_97_imag = 16'hff02;
  assign twiddle_factor_table_98_real = 16'hffdb;
  assign twiddle_factor_table_98_imag = 16'hff03;
  assign twiddle_factor_table_99_real = 16'hffcf;
  assign twiddle_factor_table_99_imag = 16'hff05;
  assign twiddle_factor_table_100_real = 16'hffc2;
  assign twiddle_factor_table_100_imag = 16'hff08;
  assign twiddle_factor_table_101_real = 16'hffb6;
  assign twiddle_factor_table_101_imag = 16'hff0c;
  assign twiddle_factor_table_102_real = 16'hffaa;
  assign twiddle_factor_table_102_imag = 16'hff0f;
  assign twiddle_factor_table_103_real = 16'hff9f;
  assign twiddle_factor_table_103_imag = 16'hff14;
  assign twiddle_factor_table_104_real = 16'hff93;
  assign twiddle_factor_table_104_imag = 16'hff19;
  assign twiddle_factor_table_105_real = 16'hff88;
  assign twiddle_factor_table_105_imag = 16'hff1f;
  assign twiddle_factor_table_106_real = 16'hff7d;
  assign twiddle_factor_table_106_imag = 16'hff25;
  assign twiddle_factor_table_107_real = 16'hff72;
  assign twiddle_factor_table_107_imag = 16'hff2c;
  assign twiddle_factor_table_108_real = 16'hff68;
  assign twiddle_factor_table_108_imag = 16'hff33;
  assign twiddle_factor_table_109_real = 16'hff5e;
  assign twiddle_factor_table_109_imag = 16'hff3b;
  assign twiddle_factor_table_110_real = 16'hff55;
  assign twiddle_factor_table_110_imag = 16'hff43;
  assign twiddle_factor_table_111_real = 16'hff4b;
  assign twiddle_factor_table_111_imag = 16'hff4b;
  assign twiddle_factor_table_112_real = 16'hff43;
  assign twiddle_factor_table_112_imag = 16'hff55;
  assign twiddle_factor_table_113_real = 16'hff3b;
  assign twiddle_factor_table_113_imag = 16'hff5e;
  assign twiddle_factor_table_114_real = 16'hff33;
  assign twiddle_factor_table_114_imag = 16'hff68;
  assign twiddle_factor_table_115_real = 16'hff2c;
  assign twiddle_factor_table_115_imag = 16'hff72;
  assign twiddle_factor_table_116_real = 16'hff25;
  assign twiddle_factor_table_116_imag = 16'hff7d;
  assign twiddle_factor_table_117_real = 16'hff1f;
  assign twiddle_factor_table_117_imag = 16'hff88;
  assign twiddle_factor_table_118_real = 16'hff19;
  assign twiddle_factor_table_118_imag = 16'hff93;
  assign twiddle_factor_table_119_real = 16'hff14;
  assign twiddle_factor_table_119_imag = 16'hff9f;
  assign twiddle_factor_table_120_real = 16'hff0f;
  assign twiddle_factor_table_120_imag = 16'hffaa;
  assign twiddle_factor_table_121_real = 16'hff0c;
  assign twiddle_factor_table_121_imag = 16'hffb6;
  assign twiddle_factor_table_122_real = 16'hff08;
  assign twiddle_factor_table_122_imag = 16'hffc2;
  assign twiddle_factor_table_123_real = 16'hff05;
  assign twiddle_factor_table_123_imag = 16'hffcf;
  assign twiddle_factor_table_124_real = 16'hff03;
  assign twiddle_factor_table_124_imag = 16'hffdb;
  assign twiddle_factor_table_125_real = 16'hff02;
  assign twiddle_factor_table_125_imag = 16'hffe7;
  assign twiddle_factor_table_126_real = 16'hff01;
  assign twiddle_factor_table_126_imag = 16'hfff4;
  assign data_reorder_0_real = data_in_0_real;
  assign data_reorder_0_imag = data_in_0_imag;
  assign data_reorder_64_real = data_in_1_real;
  assign data_reorder_64_imag = data_in_1_imag;
  assign data_reorder_32_real = data_in_2_real;
  assign data_reorder_32_imag = data_in_2_imag;
  assign data_reorder_96_real = data_in_3_real;
  assign data_reorder_96_imag = data_in_3_imag;
  assign data_reorder_16_real = data_in_4_real;
  assign data_reorder_16_imag = data_in_4_imag;
  assign data_reorder_80_real = data_in_5_real;
  assign data_reorder_80_imag = data_in_5_imag;
  assign data_reorder_48_real = data_in_6_real;
  assign data_reorder_48_imag = data_in_6_imag;
  assign data_reorder_112_real = data_in_7_real;
  assign data_reorder_112_imag = data_in_7_imag;
  assign data_reorder_8_real = data_in_8_real;
  assign data_reorder_8_imag = data_in_8_imag;
  assign data_reorder_72_real = data_in_9_real;
  assign data_reorder_72_imag = data_in_9_imag;
  assign data_reorder_40_real = data_in_10_real;
  assign data_reorder_40_imag = data_in_10_imag;
  assign data_reorder_104_real = data_in_11_real;
  assign data_reorder_104_imag = data_in_11_imag;
  assign data_reorder_24_real = data_in_12_real;
  assign data_reorder_24_imag = data_in_12_imag;
  assign data_reorder_88_real = data_in_13_real;
  assign data_reorder_88_imag = data_in_13_imag;
  assign data_reorder_56_real = data_in_14_real;
  assign data_reorder_56_imag = data_in_14_imag;
  assign data_reorder_120_real = data_in_15_real;
  assign data_reorder_120_imag = data_in_15_imag;
  assign data_reorder_4_real = data_in_16_real;
  assign data_reorder_4_imag = data_in_16_imag;
  assign data_reorder_68_real = data_in_17_real;
  assign data_reorder_68_imag = data_in_17_imag;
  assign data_reorder_36_real = data_in_18_real;
  assign data_reorder_36_imag = data_in_18_imag;
  assign data_reorder_100_real = data_in_19_real;
  assign data_reorder_100_imag = data_in_19_imag;
  assign data_reorder_20_real = data_in_20_real;
  assign data_reorder_20_imag = data_in_20_imag;
  assign data_reorder_84_real = data_in_21_real;
  assign data_reorder_84_imag = data_in_21_imag;
  assign data_reorder_52_real = data_in_22_real;
  assign data_reorder_52_imag = data_in_22_imag;
  assign data_reorder_116_real = data_in_23_real;
  assign data_reorder_116_imag = data_in_23_imag;
  assign data_reorder_12_real = data_in_24_real;
  assign data_reorder_12_imag = data_in_24_imag;
  assign data_reorder_76_real = data_in_25_real;
  assign data_reorder_76_imag = data_in_25_imag;
  assign data_reorder_44_real = data_in_26_real;
  assign data_reorder_44_imag = data_in_26_imag;
  assign data_reorder_108_real = data_in_27_real;
  assign data_reorder_108_imag = data_in_27_imag;
  assign data_reorder_28_real = data_in_28_real;
  assign data_reorder_28_imag = data_in_28_imag;
  assign data_reorder_92_real = data_in_29_real;
  assign data_reorder_92_imag = data_in_29_imag;
  assign data_reorder_60_real = data_in_30_real;
  assign data_reorder_60_imag = data_in_30_imag;
  assign data_reorder_124_real = data_in_31_real;
  assign data_reorder_124_imag = data_in_31_imag;
  assign data_reorder_2_real = data_in_32_real;
  assign data_reorder_2_imag = data_in_32_imag;
  assign data_reorder_66_real = data_in_33_real;
  assign data_reorder_66_imag = data_in_33_imag;
  assign data_reorder_34_real = data_in_34_real;
  assign data_reorder_34_imag = data_in_34_imag;
  assign data_reorder_98_real = data_in_35_real;
  assign data_reorder_98_imag = data_in_35_imag;
  assign data_reorder_18_real = data_in_36_real;
  assign data_reorder_18_imag = data_in_36_imag;
  assign data_reorder_82_real = data_in_37_real;
  assign data_reorder_82_imag = data_in_37_imag;
  assign data_reorder_50_real = data_in_38_real;
  assign data_reorder_50_imag = data_in_38_imag;
  assign data_reorder_114_real = data_in_39_real;
  assign data_reorder_114_imag = data_in_39_imag;
  assign data_reorder_10_real = data_in_40_real;
  assign data_reorder_10_imag = data_in_40_imag;
  assign data_reorder_74_real = data_in_41_real;
  assign data_reorder_74_imag = data_in_41_imag;
  assign data_reorder_42_real = data_in_42_real;
  assign data_reorder_42_imag = data_in_42_imag;
  assign data_reorder_106_real = data_in_43_real;
  assign data_reorder_106_imag = data_in_43_imag;
  assign data_reorder_26_real = data_in_44_real;
  assign data_reorder_26_imag = data_in_44_imag;
  assign data_reorder_90_real = data_in_45_real;
  assign data_reorder_90_imag = data_in_45_imag;
  assign data_reorder_58_real = data_in_46_real;
  assign data_reorder_58_imag = data_in_46_imag;
  assign data_reorder_122_real = data_in_47_real;
  assign data_reorder_122_imag = data_in_47_imag;
  assign data_reorder_6_real = data_in_48_real;
  assign data_reorder_6_imag = data_in_48_imag;
  assign data_reorder_70_real = data_in_49_real;
  assign data_reorder_70_imag = data_in_49_imag;
  assign data_reorder_38_real = data_in_50_real;
  assign data_reorder_38_imag = data_in_50_imag;
  assign data_reorder_102_real = data_in_51_real;
  assign data_reorder_102_imag = data_in_51_imag;
  assign data_reorder_22_real = data_in_52_real;
  assign data_reorder_22_imag = data_in_52_imag;
  assign data_reorder_86_real = data_in_53_real;
  assign data_reorder_86_imag = data_in_53_imag;
  assign data_reorder_54_real = data_in_54_real;
  assign data_reorder_54_imag = data_in_54_imag;
  assign data_reorder_118_real = data_in_55_real;
  assign data_reorder_118_imag = data_in_55_imag;
  assign data_reorder_14_real = data_in_56_real;
  assign data_reorder_14_imag = data_in_56_imag;
  assign data_reorder_78_real = data_in_57_real;
  assign data_reorder_78_imag = data_in_57_imag;
  assign data_reorder_46_real = data_in_58_real;
  assign data_reorder_46_imag = data_in_58_imag;
  assign data_reorder_110_real = data_in_59_real;
  assign data_reorder_110_imag = data_in_59_imag;
  assign data_reorder_30_real = data_in_60_real;
  assign data_reorder_30_imag = data_in_60_imag;
  assign data_reorder_94_real = data_in_61_real;
  assign data_reorder_94_imag = data_in_61_imag;
  assign data_reorder_62_real = data_in_62_real;
  assign data_reorder_62_imag = data_in_62_imag;
  assign data_reorder_126_real = data_in_63_real;
  assign data_reorder_126_imag = data_in_63_imag;
  assign data_reorder_1_real = data_in_64_real;
  assign data_reorder_1_imag = data_in_64_imag;
  assign data_reorder_65_real = data_in_65_real;
  assign data_reorder_65_imag = data_in_65_imag;
  assign data_reorder_33_real = data_in_66_real;
  assign data_reorder_33_imag = data_in_66_imag;
  assign data_reorder_97_real = data_in_67_real;
  assign data_reorder_97_imag = data_in_67_imag;
  assign data_reorder_17_real = data_in_68_real;
  assign data_reorder_17_imag = data_in_68_imag;
  assign data_reorder_81_real = data_in_69_real;
  assign data_reorder_81_imag = data_in_69_imag;
  assign data_reorder_49_real = data_in_70_real;
  assign data_reorder_49_imag = data_in_70_imag;
  assign data_reorder_113_real = data_in_71_real;
  assign data_reorder_113_imag = data_in_71_imag;
  assign data_reorder_9_real = data_in_72_real;
  assign data_reorder_9_imag = data_in_72_imag;
  assign data_reorder_73_real = data_in_73_real;
  assign data_reorder_73_imag = data_in_73_imag;
  assign data_reorder_41_real = data_in_74_real;
  assign data_reorder_41_imag = data_in_74_imag;
  assign data_reorder_105_real = data_in_75_real;
  assign data_reorder_105_imag = data_in_75_imag;
  assign data_reorder_25_real = data_in_76_real;
  assign data_reorder_25_imag = data_in_76_imag;
  assign data_reorder_89_real = data_in_77_real;
  assign data_reorder_89_imag = data_in_77_imag;
  assign data_reorder_57_real = data_in_78_real;
  assign data_reorder_57_imag = data_in_78_imag;
  assign data_reorder_121_real = data_in_79_real;
  assign data_reorder_121_imag = data_in_79_imag;
  assign data_reorder_5_real = data_in_80_real;
  assign data_reorder_5_imag = data_in_80_imag;
  assign data_reorder_69_real = data_in_81_real;
  assign data_reorder_69_imag = data_in_81_imag;
  assign data_reorder_37_real = data_in_82_real;
  assign data_reorder_37_imag = data_in_82_imag;
  assign data_reorder_101_real = data_in_83_real;
  assign data_reorder_101_imag = data_in_83_imag;
  assign data_reorder_21_real = data_in_84_real;
  assign data_reorder_21_imag = data_in_84_imag;
  assign data_reorder_85_real = data_in_85_real;
  assign data_reorder_85_imag = data_in_85_imag;
  assign data_reorder_53_real = data_in_86_real;
  assign data_reorder_53_imag = data_in_86_imag;
  assign data_reorder_117_real = data_in_87_real;
  assign data_reorder_117_imag = data_in_87_imag;
  assign data_reorder_13_real = data_in_88_real;
  assign data_reorder_13_imag = data_in_88_imag;
  assign data_reorder_77_real = data_in_89_real;
  assign data_reorder_77_imag = data_in_89_imag;
  assign data_reorder_45_real = data_in_90_real;
  assign data_reorder_45_imag = data_in_90_imag;
  assign data_reorder_109_real = data_in_91_real;
  assign data_reorder_109_imag = data_in_91_imag;
  assign data_reorder_29_real = data_in_92_real;
  assign data_reorder_29_imag = data_in_92_imag;
  assign data_reorder_93_real = data_in_93_real;
  assign data_reorder_93_imag = data_in_93_imag;
  assign data_reorder_61_real = data_in_94_real;
  assign data_reorder_61_imag = data_in_94_imag;
  assign data_reorder_125_real = data_in_95_real;
  assign data_reorder_125_imag = data_in_95_imag;
  assign data_reorder_3_real = data_in_96_real;
  assign data_reorder_3_imag = data_in_96_imag;
  assign data_reorder_67_real = data_in_97_real;
  assign data_reorder_67_imag = data_in_97_imag;
  assign data_reorder_35_real = data_in_98_real;
  assign data_reorder_35_imag = data_in_98_imag;
  assign data_reorder_99_real = data_in_99_real;
  assign data_reorder_99_imag = data_in_99_imag;
  assign data_reorder_19_real = data_in_100_real;
  assign data_reorder_19_imag = data_in_100_imag;
  assign data_reorder_83_real = data_in_101_real;
  assign data_reorder_83_imag = data_in_101_imag;
  assign data_reorder_51_real = data_in_102_real;
  assign data_reorder_51_imag = data_in_102_imag;
  assign data_reorder_115_real = data_in_103_real;
  assign data_reorder_115_imag = data_in_103_imag;
  assign data_reorder_11_real = data_in_104_real;
  assign data_reorder_11_imag = data_in_104_imag;
  assign data_reorder_75_real = data_in_105_real;
  assign data_reorder_75_imag = data_in_105_imag;
  assign data_reorder_43_real = data_in_106_real;
  assign data_reorder_43_imag = data_in_106_imag;
  assign data_reorder_107_real = data_in_107_real;
  assign data_reorder_107_imag = data_in_107_imag;
  assign data_reorder_27_real = data_in_108_real;
  assign data_reorder_27_imag = data_in_108_imag;
  assign data_reorder_91_real = data_in_109_real;
  assign data_reorder_91_imag = data_in_109_imag;
  assign data_reorder_59_real = data_in_110_real;
  assign data_reorder_59_imag = data_in_110_imag;
  assign data_reorder_123_real = data_in_111_real;
  assign data_reorder_123_imag = data_in_111_imag;
  assign data_reorder_7_real = data_in_112_real;
  assign data_reorder_7_imag = data_in_112_imag;
  assign data_reorder_71_real = data_in_113_real;
  assign data_reorder_71_imag = data_in_113_imag;
  assign data_reorder_39_real = data_in_114_real;
  assign data_reorder_39_imag = data_in_114_imag;
  assign data_reorder_103_real = data_in_115_real;
  assign data_reorder_103_imag = data_in_115_imag;
  assign data_reorder_23_real = data_in_116_real;
  assign data_reorder_23_imag = data_in_116_imag;
  assign data_reorder_87_real = data_in_117_real;
  assign data_reorder_87_imag = data_in_117_imag;
  assign data_reorder_55_real = data_in_118_real;
  assign data_reorder_55_imag = data_in_118_imag;
  assign data_reorder_119_real = data_in_119_real;
  assign data_reorder_119_imag = data_in_119_imag;
  assign data_reorder_15_real = data_in_120_real;
  assign data_reorder_15_imag = data_in_120_imag;
  assign data_reorder_79_real = data_in_121_real;
  assign data_reorder_79_imag = data_in_121_imag;
  assign data_reorder_47_real = data_in_122_real;
  assign data_reorder_47_imag = data_in_122_imag;
  assign data_reorder_111_real = data_in_123_real;
  assign data_reorder_111_imag = data_in_123_imag;
  assign data_reorder_31_real = data_in_124_real;
  assign data_reorder_31_imag = data_in_124_imag;
  assign data_reorder_95_real = data_in_125_real;
  assign data_reorder_95_imag = data_in_125_imag;
  assign data_reorder_63_real = data_in_126_real;
  assign data_reorder_63_imag = data_in_126_imag;
  assign data_reorder_127_real = data_in_127_real;
  assign data_reorder_127_imag = data_in_127_imag;
  always @ (*) begin
    current_level_cnt_willIncrement = 1'b0;
    if(current_level_cond_period)begin
      current_level_cnt_willIncrement = 1'b1;
    end
  end

  assign current_level_cnt_willClear = 1'b0;
  assign current_level_cnt_willOverflowIfInc = (current_level_cnt_value == 3'b111);
  assign current_level_cnt_willOverflow = (current_level_cnt_willOverflowIfInc && current_level_cnt_willIncrement);
  always @ (*) begin
    current_level_cnt_valueNext = (current_level_cnt_value + _zz_2690);
    if(current_level_cnt_willClear)begin
      current_level_cnt_valueNext = 3'b000;
    end
  end

  assign current_level_cond_period = (io_data_in_valid_regNext || current_level_cond_period_minus_1);
  assign _zz_1793 = ($signed(_zz_2691) - $signed(_zz_2692));
  assign _zz_1 = _zz_2693[15 : 0];
  assign _zz_1794 = ($signed(_zz_2694) + $signed(_zz_2695));
  assign _zz_2 = _zz_2696[15 : 0];
  assign _zz_3 = 1'b1;
  assign _zz_4 = 1'b1;
  assign _zz_1795 = ($signed(_zz_2713) - $signed(_zz_2714));
  assign _zz_5 = _zz_2715[15 : 0];
  assign _zz_1796 = ($signed(_zz_2716) + $signed(_zz_2717));
  assign _zz_6 = _zz_2718[15 : 0];
  assign _zz_7 = 1'b1;
  assign _zz_8 = 1'b1;
  assign _zz_1797 = ($signed(_zz_2735) - $signed(_zz_2736));
  assign _zz_9 = _zz_2737[15 : 0];
  assign _zz_1798 = ($signed(_zz_2738) + $signed(_zz_2739));
  assign _zz_10 = _zz_2740[15 : 0];
  assign _zz_11 = 1'b1;
  assign _zz_12 = 1'b1;
  assign _zz_1799 = ($signed(_zz_2757) - $signed(_zz_2758));
  assign _zz_13 = _zz_2759[15 : 0];
  assign _zz_1800 = ($signed(_zz_2760) + $signed(_zz_2761));
  assign _zz_14 = _zz_2762[15 : 0];
  assign _zz_15 = 1'b1;
  assign _zz_16 = 1'b1;
  assign _zz_1801 = ($signed(_zz_2779) - $signed(_zz_2780));
  assign _zz_17 = _zz_2781[15 : 0];
  assign _zz_1802 = ($signed(_zz_2782) + $signed(_zz_2783));
  assign _zz_18 = _zz_2784[15 : 0];
  assign _zz_19 = 1'b1;
  assign _zz_20 = 1'b1;
  assign _zz_1803 = ($signed(_zz_2801) - $signed(_zz_2802));
  assign _zz_21 = _zz_2803[15 : 0];
  assign _zz_1804 = ($signed(_zz_2804) + $signed(_zz_2805));
  assign _zz_22 = _zz_2806[15 : 0];
  assign _zz_23 = 1'b1;
  assign _zz_24 = 1'b1;
  assign _zz_1805 = ($signed(_zz_2823) - $signed(_zz_2824));
  assign _zz_25 = _zz_2825[15 : 0];
  assign _zz_1806 = ($signed(_zz_2826) + $signed(_zz_2827));
  assign _zz_26 = _zz_2828[15 : 0];
  assign _zz_27 = 1'b1;
  assign _zz_28 = 1'b1;
  assign _zz_1807 = ($signed(_zz_2845) - $signed(_zz_2846));
  assign _zz_29 = _zz_2847[15 : 0];
  assign _zz_1808 = ($signed(_zz_2848) + $signed(_zz_2849));
  assign _zz_30 = _zz_2850[15 : 0];
  assign _zz_31 = 1'b1;
  assign _zz_32 = 1'b1;
  assign _zz_1809 = ($signed(_zz_2867) - $signed(_zz_2868));
  assign _zz_33 = _zz_2869[15 : 0];
  assign _zz_1810 = ($signed(_zz_2870) + $signed(_zz_2871));
  assign _zz_34 = _zz_2872[15 : 0];
  assign _zz_35 = 1'b1;
  assign _zz_36 = 1'b1;
  assign _zz_1811 = ($signed(_zz_2889) - $signed(_zz_2890));
  assign _zz_37 = _zz_2891[15 : 0];
  assign _zz_1812 = ($signed(_zz_2892) + $signed(_zz_2893));
  assign _zz_38 = _zz_2894[15 : 0];
  assign _zz_39 = 1'b1;
  assign _zz_40 = 1'b1;
  assign _zz_1813 = ($signed(_zz_2911) - $signed(_zz_2912));
  assign _zz_41 = _zz_2913[15 : 0];
  assign _zz_1814 = ($signed(_zz_2914) + $signed(_zz_2915));
  assign _zz_42 = _zz_2916[15 : 0];
  assign _zz_43 = 1'b1;
  assign _zz_44 = 1'b1;
  assign _zz_1815 = ($signed(_zz_2933) - $signed(_zz_2934));
  assign _zz_45 = _zz_2935[15 : 0];
  assign _zz_1816 = ($signed(_zz_2936) + $signed(_zz_2937));
  assign _zz_46 = _zz_2938[15 : 0];
  assign _zz_47 = 1'b1;
  assign _zz_48 = 1'b1;
  assign _zz_1817 = ($signed(_zz_2955) - $signed(_zz_2956));
  assign _zz_49 = _zz_2957[15 : 0];
  assign _zz_1818 = ($signed(_zz_2958) + $signed(_zz_2959));
  assign _zz_50 = _zz_2960[15 : 0];
  assign _zz_51 = 1'b1;
  assign _zz_52 = 1'b1;
  assign _zz_1819 = ($signed(_zz_2977) - $signed(_zz_2978));
  assign _zz_53 = _zz_2979[15 : 0];
  assign _zz_1820 = ($signed(_zz_2980) + $signed(_zz_2981));
  assign _zz_54 = _zz_2982[15 : 0];
  assign _zz_55 = 1'b1;
  assign _zz_56 = 1'b1;
  assign _zz_1821 = ($signed(_zz_2999) - $signed(_zz_3000));
  assign _zz_57 = _zz_3001[15 : 0];
  assign _zz_1822 = ($signed(_zz_3002) + $signed(_zz_3003));
  assign _zz_58 = _zz_3004[15 : 0];
  assign _zz_59 = 1'b1;
  assign _zz_60 = 1'b1;
  assign _zz_1823 = ($signed(_zz_3021) - $signed(_zz_3022));
  assign _zz_61 = _zz_3023[15 : 0];
  assign _zz_1824 = ($signed(_zz_3024) + $signed(_zz_3025));
  assign _zz_62 = _zz_3026[15 : 0];
  assign _zz_63 = 1'b1;
  assign _zz_64 = 1'b1;
  assign _zz_1825 = ($signed(_zz_3043) - $signed(_zz_3044));
  assign _zz_65 = _zz_3045[15 : 0];
  assign _zz_1826 = ($signed(_zz_3046) + $signed(_zz_3047));
  assign _zz_66 = _zz_3048[15 : 0];
  assign _zz_67 = 1'b1;
  assign _zz_68 = 1'b1;
  assign _zz_1827 = ($signed(_zz_3065) - $signed(_zz_3066));
  assign _zz_69 = _zz_3067[15 : 0];
  assign _zz_1828 = ($signed(_zz_3068) + $signed(_zz_3069));
  assign _zz_70 = _zz_3070[15 : 0];
  assign _zz_71 = 1'b1;
  assign _zz_72 = 1'b1;
  assign _zz_1829 = ($signed(_zz_3087) - $signed(_zz_3088));
  assign _zz_73 = _zz_3089[15 : 0];
  assign _zz_1830 = ($signed(_zz_3090) + $signed(_zz_3091));
  assign _zz_74 = _zz_3092[15 : 0];
  assign _zz_75 = 1'b1;
  assign _zz_76 = 1'b1;
  assign _zz_1831 = ($signed(_zz_3109) - $signed(_zz_3110));
  assign _zz_77 = _zz_3111[15 : 0];
  assign _zz_1832 = ($signed(_zz_3112) + $signed(_zz_3113));
  assign _zz_78 = _zz_3114[15 : 0];
  assign _zz_79 = 1'b1;
  assign _zz_80 = 1'b1;
  assign _zz_1833 = ($signed(_zz_3131) - $signed(_zz_3132));
  assign _zz_81 = _zz_3133[15 : 0];
  assign _zz_1834 = ($signed(_zz_3134) + $signed(_zz_3135));
  assign _zz_82 = _zz_3136[15 : 0];
  assign _zz_83 = 1'b1;
  assign _zz_84 = 1'b1;
  assign _zz_1835 = ($signed(_zz_3153) - $signed(_zz_3154));
  assign _zz_85 = _zz_3155[15 : 0];
  assign _zz_1836 = ($signed(_zz_3156) + $signed(_zz_3157));
  assign _zz_86 = _zz_3158[15 : 0];
  assign _zz_87 = 1'b1;
  assign _zz_88 = 1'b1;
  assign _zz_1837 = ($signed(_zz_3175) - $signed(_zz_3176));
  assign _zz_89 = _zz_3177[15 : 0];
  assign _zz_1838 = ($signed(_zz_3178) + $signed(_zz_3179));
  assign _zz_90 = _zz_3180[15 : 0];
  assign _zz_91 = 1'b1;
  assign _zz_92 = 1'b1;
  assign _zz_1839 = ($signed(_zz_3197) - $signed(_zz_3198));
  assign _zz_93 = _zz_3199[15 : 0];
  assign _zz_1840 = ($signed(_zz_3200) + $signed(_zz_3201));
  assign _zz_94 = _zz_3202[15 : 0];
  assign _zz_95 = 1'b1;
  assign _zz_96 = 1'b1;
  assign _zz_1841 = ($signed(_zz_3219) - $signed(_zz_3220));
  assign _zz_97 = _zz_3221[15 : 0];
  assign _zz_1842 = ($signed(_zz_3222) + $signed(_zz_3223));
  assign _zz_98 = _zz_3224[15 : 0];
  assign _zz_99 = 1'b1;
  assign _zz_100 = 1'b1;
  assign _zz_1843 = ($signed(_zz_3241) - $signed(_zz_3242));
  assign _zz_101 = _zz_3243[15 : 0];
  assign _zz_1844 = ($signed(_zz_3244) + $signed(_zz_3245));
  assign _zz_102 = _zz_3246[15 : 0];
  assign _zz_103 = 1'b1;
  assign _zz_104 = 1'b1;
  assign _zz_1845 = ($signed(_zz_3263) - $signed(_zz_3264));
  assign _zz_105 = _zz_3265[15 : 0];
  assign _zz_1846 = ($signed(_zz_3266) + $signed(_zz_3267));
  assign _zz_106 = _zz_3268[15 : 0];
  assign _zz_107 = 1'b1;
  assign _zz_108 = 1'b1;
  assign _zz_1847 = ($signed(_zz_3285) - $signed(_zz_3286));
  assign _zz_109 = _zz_3287[15 : 0];
  assign _zz_1848 = ($signed(_zz_3288) + $signed(_zz_3289));
  assign _zz_110 = _zz_3290[15 : 0];
  assign _zz_111 = 1'b1;
  assign _zz_112 = 1'b1;
  assign _zz_1849 = ($signed(_zz_3307) - $signed(_zz_3308));
  assign _zz_113 = _zz_3309[15 : 0];
  assign _zz_1850 = ($signed(_zz_3310) + $signed(_zz_3311));
  assign _zz_114 = _zz_3312[15 : 0];
  assign _zz_115 = 1'b1;
  assign _zz_116 = 1'b1;
  assign _zz_1851 = ($signed(_zz_3329) - $signed(_zz_3330));
  assign _zz_117 = _zz_3331[15 : 0];
  assign _zz_1852 = ($signed(_zz_3332) + $signed(_zz_3333));
  assign _zz_118 = _zz_3334[15 : 0];
  assign _zz_119 = 1'b1;
  assign _zz_120 = 1'b1;
  assign _zz_1853 = ($signed(_zz_3351) - $signed(_zz_3352));
  assign _zz_121 = _zz_3353[15 : 0];
  assign _zz_1854 = ($signed(_zz_3354) + $signed(_zz_3355));
  assign _zz_122 = _zz_3356[15 : 0];
  assign _zz_123 = 1'b1;
  assign _zz_124 = 1'b1;
  assign _zz_1855 = ($signed(_zz_3373) - $signed(_zz_3374));
  assign _zz_125 = _zz_3375[15 : 0];
  assign _zz_1856 = ($signed(_zz_3376) + $signed(_zz_3377));
  assign _zz_126 = _zz_3378[15 : 0];
  assign _zz_127 = 1'b1;
  assign _zz_128 = 1'b1;
  assign _zz_1857 = ($signed(_zz_3395) - $signed(_zz_3396));
  assign _zz_129 = _zz_3397[15 : 0];
  assign _zz_1858 = ($signed(_zz_3398) + $signed(_zz_3399));
  assign _zz_130 = _zz_3400[15 : 0];
  assign _zz_131 = 1'b1;
  assign _zz_132 = 1'b1;
  assign _zz_1859 = ($signed(_zz_3417) - $signed(_zz_3418));
  assign _zz_133 = _zz_3419[15 : 0];
  assign _zz_1860 = ($signed(_zz_3420) + $signed(_zz_3421));
  assign _zz_134 = _zz_3422[15 : 0];
  assign _zz_135 = 1'b1;
  assign _zz_136 = 1'b1;
  assign _zz_1861 = ($signed(_zz_3439) - $signed(_zz_3440));
  assign _zz_137 = _zz_3441[15 : 0];
  assign _zz_1862 = ($signed(_zz_3442) + $signed(_zz_3443));
  assign _zz_138 = _zz_3444[15 : 0];
  assign _zz_139 = 1'b1;
  assign _zz_140 = 1'b1;
  assign _zz_1863 = ($signed(_zz_3461) - $signed(_zz_3462));
  assign _zz_141 = _zz_3463[15 : 0];
  assign _zz_1864 = ($signed(_zz_3464) + $signed(_zz_3465));
  assign _zz_142 = _zz_3466[15 : 0];
  assign _zz_143 = 1'b1;
  assign _zz_144 = 1'b1;
  assign _zz_1865 = ($signed(_zz_3483) - $signed(_zz_3484));
  assign _zz_145 = _zz_3485[15 : 0];
  assign _zz_1866 = ($signed(_zz_3486) + $signed(_zz_3487));
  assign _zz_146 = _zz_3488[15 : 0];
  assign _zz_147 = 1'b1;
  assign _zz_148 = 1'b1;
  assign _zz_1867 = ($signed(_zz_3505) - $signed(_zz_3506));
  assign _zz_149 = _zz_3507[15 : 0];
  assign _zz_1868 = ($signed(_zz_3508) + $signed(_zz_3509));
  assign _zz_150 = _zz_3510[15 : 0];
  assign _zz_151 = 1'b1;
  assign _zz_152 = 1'b1;
  assign _zz_1869 = ($signed(_zz_3527) - $signed(_zz_3528));
  assign _zz_153 = _zz_3529[15 : 0];
  assign _zz_1870 = ($signed(_zz_3530) + $signed(_zz_3531));
  assign _zz_154 = _zz_3532[15 : 0];
  assign _zz_155 = 1'b1;
  assign _zz_156 = 1'b1;
  assign _zz_1871 = ($signed(_zz_3549) - $signed(_zz_3550));
  assign _zz_157 = _zz_3551[15 : 0];
  assign _zz_1872 = ($signed(_zz_3552) + $signed(_zz_3553));
  assign _zz_158 = _zz_3554[15 : 0];
  assign _zz_159 = 1'b1;
  assign _zz_160 = 1'b1;
  assign _zz_1873 = ($signed(_zz_3571) - $signed(_zz_3572));
  assign _zz_161 = _zz_3573[15 : 0];
  assign _zz_1874 = ($signed(_zz_3574) + $signed(_zz_3575));
  assign _zz_162 = _zz_3576[15 : 0];
  assign _zz_163 = 1'b1;
  assign _zz_164 = 1'b1;
  assign _zz_1875 = ($signed(_zz_3593) - $signed(_zz_3594));
  assign _zz_165 = _zz_3595[15 : 0];
  assign _zz_1876 = ($signed(_zz_3596) + $signed(_zz_3597));
  assign _zz_166 = _zz_3598[15 : 0];
  assign _zz_167 = 1'b1;
  assign _zz_168 = 1'b1;
  assign _zz_1877 = ($signed(_zz_3615) - $signed(_zz_3616));
  assign _zz_169 = _zz_3617[15 : 0];
  assign _zz_1878 = ($signed(_zz_3618) + $signed(_zz_3619));
  assign _zz_170 = _zz_3620[15 : 0];
  assign _zz_171 = 1'b1;
  assign _zz_172 = 1'b1;
  assign _zz_1879 = ($signed(_zz_3637) - $signed(_zz_3638));
  assign _zz_173 = _zz_3639[15 : 0];
  assign _zz_1880 = ($signed(_zz_3640) + $signed(_zz_3641));
  assign _zz_174 = _zz_3642[15 : 0];
  assign _zz_175 = 1'b1;
  assign _zz_176 = 1'b1;
  assign _zz_1881 = ($signed(_zz_3659) - $signed(_zz_3660));
  assign _zz_177 = _zz_3661[15 : 0];
  assign _zz_1882 = ($signed(_zz_3662) + $signed(_zz_3663));
  assign _zz_178 = _zz_3664[15 : 0];
  assign _zz_179 = 1'b1;
  assign _zz_180 = 1'b1;
  assign _zz_1883 = ($signed(_zz_3681) - $signed(_zz_3682));
  assign _zz_181 = _zz_3683[15 : 0];
  assign _zz_1884 = ($signed(_zz_3684) + $signed(_zz_3685));
  assign _zz_182 = _zz_3686[15 : 0];
  assign _zz_183 = 1'b1;
  assign _zz_184 = 1'b1;
  assign _zz_1885 = ($signed(_zz_3703) - $signed(_zz_3704));
  assign _zz_185 = _zz_3705[15 : 0];
  assign _zz_1886 = ($signed(_zz_3706) + $signed(_zz_3707));
  assign _zz_186 = _zz_3708[15 : 0];
  assign _zz_187 = 1'b1;
  assign _zz_188 = 1'b1;
  assign _zz_1887 = ($signed(_zz_3725) - $signed(_zz_3726));
  assign _zz_189 = _zz_3727[15 : 0];
  assign _zz_1888 = ($signed(_zz_3728) + $signed(_zz_3729));
  assign _zz_190 = _zz_3730[15 : 0];
  assign _zz_191 = 1'b1;
  assign _zz_192 = 1'b1;
  assign _zz_1889 = ($signed(_zz_3747) - $signed(_zz_3748));
  assign _zz_193 = _zz_3749[15 : 0];
  assign _zz_1890 = ($signed(_zz_3750) + $signed(_zz_3751));
  assign _zz_194 = _zz_3752[15 : 0];
  assign _zz_195 = 1'b1;
  assign _zz_196 = 1'b1;
  assign _zz_1891 = ($signed(_zz_3769) - $signed(_zz_3770));
  assign _zz_197 = _zz_3771[15 : 0];
  assign _zz_1892 = ($signed(_zz_3772) + $signed(_zz_3773));
  assign _zz_198 = _zz_3774[15 : 0];
  assign _zz_199 = 1'b1;
  assign _zz_200 = 1'b1;
  assign _zz_1893 = ($signed(_zz_3791) - $signed(_zz_3792));
  assign _zz_201 = _zz_3793[15 : 0];
  assign _zz_1894 = ($signed(_zz_3794) + $signed(_zz_3795));
  assign _zz_202 = _zz_3796[15 : 0];
  assign _zz_203 = 1'b1;
  assign _zz_204 = 1'b1;
  assign _zz_1895 = ($signed(_zz_3813) - $signed(_zz_3814));
  assign _zz_205 = _zz_3815[15 : 0];
  assign _zz_1896 = ($signed(_zz_3816) + $signed(_zz_3817));
  assign _zz_206 = _zz_3818[15 : 0];
  assign _zz_207 = 1'b1;
  assign _zz_208 = 1'b1;
  assign _zz_1897 = ($signed(_zz_3835) - $signed(_zz_3836));
  assign _zz_209 = _zz_3837[15 : 0];
  assign _zz_1898 = ($signed(_zz_3838) + $signed(_zz_3839));
  assign _zz_210 = _zz_3840[15 : 0];
  assign _zz_211 = 1'b1;
  assign _zz_212 = 1'b1;
  assign _zz_1899 = ($signed(_zz_3857) - $signed(_zz_3858));
  assign _zz_213 = _zz_3859[15 : 0];
  assign _zz_1900 = ($signed(_zz_3860) + $signed(_zz_3861));
  assign _zz_214 = _zz_3862[15 : 0];
  assign _zz_215 = 1'b1;
  assign _zz_216 = 1'b1;
  assign _zz_1901 = ($signed(_zz_3879) - $signed(_zz_3880));
  assign _zz_217 = _zz_3881[15 : 0];
  assign _zz_1902 = ($signed(_zz_3882) + $signed(_zz_3883));
  assign _zz_218 = _zz_3884[15 : 0];
  assign _zz_219 = 1'b1;
  assign _zz_220 = 1'b1;
  assign _zz_1903 = ($signed(_zz_3901) - $signed(_zz_3902));
  assign _zz_221 = _zz_3903[15 : 0];
  assign _zz_1904 = ($signed(_zz_3904) + $signed(_zz_3905));
  assign _zz_222 = _zz_3906[15 : 0];
  assign _zz_223 = 1'b1;
  assign _zz_224 = 1'b1;
  assign _zz_1905 = ($signed(_zz_3923) - $signed(_zz_3924));
  assign _zz_225 = _zz_3925[15 : 0];
  assign _zz_1906 = ($signed(_zz_3926) + $signed(_zz_3927));
  assign _zz_226 = _zz_3928[15 : 0];
  assign _zz_227 = 1'b1;
  assign _zz_228 = 1'b1;
  assign _zz_1907 = ($signed(_zz_3945) - $signed(_zz_3946));
  assign _zz_229 = _zz_3947[15 : 0];
  assign _zz_1908 = ($signed(_zz_3948) + $signed(_zz_3949));
  assign _zz_230 = _zz_3950[15 : 0];
  assign _zz_231 = 1'b1;
  assign _zz_232 = 1'b1;
  assign _zz_1909 = ($signed(_zz_3967) - $signed(_zz_3968));
  assign _zz_233 = _zz_3969[15 : 0];
  assign _zz_1910 = ($signed(_zz_3970) + $signed(_zz_3971));
  assign _zz_234 = _zz_3972[15 : 0];
  assign _zz_235 = 1'b1;
  assign _zz_236 = 1'b1;
  assign _zz_1911 = ($signed(_zz_3989) - $signed(_zz_3990));
  assign _zz_237 = _zz_3991[15 : 0];
  assign _zz_1912 = ($signed(_zz_3992) + $signed(_zz_3993));
  assign _zz_238 = _zz_3994[15 : 0];
  assign _zz_239 = 1'b1;
  assign _zz_240 = 1'b1;
  assign _zz_1913 = ($signed(_zz_4011) - $signed(_zz_4012));
  assign _zz_241 = _zz_4013[15 : 0];
  assign _zz_1914 = ($signed(_zz_4014) + $signed(_zz_4015));
  assign _zz_242 = _zz_4016[15 : 0];
  assign _zz_243 = 1'b1;
  assign _zz_244 = 1'b1;
  assign _zz_1915 = ($signed(_zz_4033) - $signed(_zz_4034));
  assign _zz_245 = _zz_4035[15 : 0];
  assign _zz_1916 = ($signed(_zz_4036) + $signed(_zz_4037));
  assign _zz_246 = _zz_4038[15 : 0];
  assign _zz_247 = 1'b1;
  assign _zz_248 = 1'b1;
  assign _zz_1917 = ($signed(_zz_4055) - $signed(_zz_4056));
  assign _zz_249 = _zz_4057[15 : 0];
  assign _zz_1918 = ($signed(_zz_4058) + $signed(_zz_4059));
  assign _zz_250 = _zz_4060[15 : 0];
  assign _zz_251 = 1'b1;
  assign _zz_252 = 1'b1;
  assign _zz_1919 = ($signed(_zz_4077) - $signed(_zz_4078));
  assign _zz_253 = _zz_4079[15 : 0];
  assign _zz_1920 = ($signed(_zz_4080) + $signed(_zz_4081));
  assign _zz_254 = _zz_4082[15 : 0];
  assign _zz_255 = 1'b1;
  assign _zz_256 = 1'b1;
  assign _zz_1921 = ($signed(_zz_4099) - $signed(_zz_4100));
  assign _zz_257 = _zz_4101[15 : 0];
  assign _zz_1922 = ($signed(_zz_4102) + $signed(_zz_4103));
  assign _zz_258 = _zz_4104[15 : 0];
  assign _zz_259 = 1'b1;
  assign _zz_260 = 1'b1;
  assign _zz_1923 = ($signed(_zz_4121) - $signed(_zz_4122));
  assign _zz_261 = _zz_4123[15 : 0];
  assign _zz_1924 = ($signed(_zz_4124) + $signed(_zz_4125));
  assign _zz_262 = _zz_4126[15 : 0];
  assign _zz_263 = 1'b1;
  assign _zz_264 = 1'b1;
  assign _zz_1925 = ($signed(_zz_4143) - $signed(_zz_4144));
  assign _zz_265 = _zz_4145[15 : 0];
  assign _zz_1926 = ($signed(_zz_4146) + $signed(_zz_4147));
  assign _zz_266 = _zz_4148[15 : 0];
  assign _zz_267 = 1'b1;
  assign _zz_268 = 1'b1;
  assign _zz_1927 = ($signed(_zz_4165) - $signed(_zz_4166));
  assign _zz_269 = _zz_4167[15 : 0];
  assign _zz_1928 = ($signed(_zz_4168) + $signed(_zz_4169));
  assign _zz_270 = _zz_4170[15 : 0];
  assign _zz_271 = 1'b1;
  assign _zz_272 = 1'b1;
  assign _zz_1929 = ($signed(_zz_4187) - $signed(_zz_4188));
  assign _zz_273 = _zz_4189[15 : 0];
  assign _zz_1930 = ($signed(_zz_4190) + $signed(_zz_4191));
  assign _zz_274 = _zz_4192[15 : 0];
  assign _zz_275 = 1'b1;
  assign _zz_276 = 1'b1;
  assign _zz_1931 = ($signed(_zz_4209) - $signed(_zz_4210));
  assign _zz_277 = _zz_4211[15 : 0];
  assign _zz_1932 = ($signed(_zz_4212) + $signed(_zz_4213));
  assign _zz_278 = _zz_4214[15 : 0];
  assign _zz_279 = 1'b1;
  assign _zz_280 = 1'b1;
  assign _zz_1933 = ($signed(_zz_4231) - $signed(_zz_4232));
  assign _zz_281 = _zz_4233[15 : 0];
  assign _zz_1934 = ($signed(_zz_4234) + $signed(_zz_4235));
  assign _zz_282 = _zz_4236[15 : 0];
  assign _zz_283 = 1'b1;
  assign _zz_284 = 1'b1;
  assign _zz_1935 = ($signed(_zz_4253) - $signed(_zz_4254));
  assign _zz_285 = _zz_4255[15 : 0];
  assign _zz_1936 = ($signed(_zz_4256) + $signed(_zz_4257));
  assign _zz_286 = _zz_4258[15 : 0];
  assign _zz_287 = 1'b1;
  assign _zz_288 = 1'b1;
  assign _zz_1937 = ($signed(_zz_4275) - $signed(_zz_4276));
  assign _zz_289 = _zz_4277[15 : 0];
  assign _zz_1938 = ($signed(_zz_4278) + $signed(_zz_4279));
  assign _zz_290 = _zz_4280[15 : 0];
  assign _zz_291 = 1'b1;
  assign _zz_292 = 1'b1;
  assign _zz_1939 = ($signed(_zz_4297) - $signed(_zz_4298));
  assign _zz_293 = _zz_4299[15 : 0];
  assign _zz_1940 = ($signed(_zz_4300) + $signed(_zz_4301));
  assign _zz_294 = _zz_4302[15 : 0];
  assign _zz_295 = 1'b1;
  assign _zz_296 = 1'b1;
  assign _zz_1941 = ($signed(_zz_4319) - $signed(_zz_4320));
  assign _zz_297 = _zz_4321[15 : 0];
  assign _zz_1942 = ($signed(_zz_4322) + $signed(_zz_4323));
  assign _zz_298 = _zz_4324[15 : 0];
  assign _zz_299 = 1'b1;
  assign _zz_300 = 1'b1;
  assign _zz_1943 = ($signed(_zz_4341) - $signed(_zz_4342));
  assign _zz_301 = _zz_4343[15 : 0];
  assign _zz_1944 = ($signed(_zz_4344) + $signed(_zz_4345));
  assign _zz_302 = _zz_4346[15 : 0];
  assign _zz_303 = 1'b1;
  assign _zz_304 = 1'b1;
  assign _zz_1945 = ($signed(_zz_4363) - $signed(_zz_4364));
  assign _zz_305 = _zz_4365[15 : 0];
  assign _zz_1946 = ($signed(_zz_4366) + $signed(_zz_4367));
  assign _zz_306 = _zz_4368[15 : 0];
  assign _zz_307 = 1'b1;
  assign _zz_308 = 1'b1;
  assign _zz_1947 = ($signed(_zz_4385) - $signed(_zz_4386));
  assign _zz_309 = _zz_4387[15 : 0];
  assign _zz_1948 = ($signed(_zz_4388) + $signed(_zz_4389));
  assign _zz_310 = _zz_4390[15 : 0];
  assign _zz_311 = 1'b1;
  assign _zz_312 = 1'b1;
  assign _zz_1949 = ($signed(_zz_4407) - $signed(_zz_4408));
  assign _zz_313 = _zz_4409[15 : 0];
  assign _zz_1950 = ($signed(_zz_4410) + $signed(_zz_4411));
  assign _zz_314 = _zz_4412[15 : 0];
  assign _zz_315 = 1'b1;
  assign _zz_316 = 1'b1;
  assign _zz_1951 = ($signed(_zz_4429) - $signed(_zz_4430));
  assign _zz_317 = _zz_4431[15 : 0];
  assign _zz_1952 = ($signed(_zz_4432) + $signed(_zz_4433));
  assign _zz_318 = _zz_4434[15 : 0];
  assign _zz_319 = 1'b1;
  assign _zz_320 = 1'b1;
  assign _zz_1953 = ($signed(_zz_4451) - $signed(_zz_4452));
  assign _zz_321 = _zz_4453[15 : 0];
  assign _zz_1954 = ($signed(_zz_4454) + $signed(_zz_4455));
  assign _zz_322 = _zz_4456[15 : 0];
  assign _zz_323 = 1'b1;
  assign _zz_324 = 1'b1;
  assign _zz_1955 = ($signed(_zz_4473) - $signed(_zz_4474));
  assign _zz_325 = _zz_4475[15 : 0];
  assign _zz_1956 = ($signed(_zz_4476) + $signed(_zz_4477));
  assign _zz_326 = _zz_4478[15 : 0];
  assign _zz_327 = 1'b1;
  assign _zz_328 = 1'b1;
  assign _zz_1957 = ($signed(_zz_4495) - $signed(_zz_4496));
  assign _zz_329 = _zz_4497[15 : 0];
  assign _zz_1958 = ($signed(_zz_4498) + $signed(_zz_4499));
  assign _zz_330 = _zz_4500[15 : 0];
  assign _zz_331 = 1'b1;
  assign _zz_332 = 1'b1;
  assign _zz_1959 = ($signed(_zz_4517) - $signed(_zz_4518));
  assign _zz_333 = _zz_4519[15 : 0];
  assign _zz_1960 = ($signed(_zz_4520) + $signed(_zz_4521));
  assign _zz_334 = _zz_4522[15 : 0];
  assign _zz_335 = 1'b1;
  assign _zz_336 = 1'b1;
  assign _zz_1961 = ($signed(_zz_4539) - $signed(_zz_4540));
  assign _zz_337 = _zz_4541[15 : 0];
  assign _zz_1962 = ($signed(_zz_4542) + $signed(_zz_4543));
  assign _zz_338 = _zz_4544[15 : 0];
  assign _zz_339 = 1'b1;
  assign _zz_340 = 1'b1;
  assign _zz_1963 = ($signed(_zz_4561) - $signed(_zz_4562));
  assign _zz_341 = _zz_4563[15 : 0];
  assign _zz_1964 = ($signed(_zz_4564) + $signed(_zz_4565));
  assign _zz_342 = _zz_4566[15 : 0];
  assign _zz_343 = 1'b1;
  assign _zz_344 = 1'b1;
  assign _zz_1965 = ($signed(_zz_4583) - $signed(_zz_4584));
  assign _zz_345 = _zz_4585[15 : 0];
  assign _zz_1966 = ($signed(_zz_4586) + $signed(_zz_4587));
  assign _zz_346 = _zz_4588[15 : 0];
  assign _zz_347 = 1'b1;
  assign _zz_348 = 1'b1;
  assign _zz_1967 = ($signed(_zz_4605) - $signed(_zz_4606));
  assign _zz_349 = _zz_4607[15 : 0];
  assign _zz_1968 = ($signed(_zz_4608) + $signed(_zz_4609));
  assign _zz_350 = _zz_4610[15 : 0];
  assign _zz_351 = 1'b1;
  assign _zz_352 = 1'b1;
  assign _zz_1969 = ($signed(_zz_4627) - $signed(_zz_4628));
  assign _zz_353 = _zz_4629[15 : 0];
  assign _zz_1970 = ($signed(_zz_4630) + $signed(_zz_4631));
  assign _zz_354 = _zz_4632[15 : 0];
  assign _zz_355 = 1'b1;
  assign _zz_356 = 1'b1;
  assign _zz_1971 = ($signed(_zz_4649) - $signed(_zz_4650));
  assign _zz_357 = _zz_4651[15 : 0];
  assign _zz_1972 = ($signed(_zz_4652) + $signed(_zz_4653));
  assign _zz_358 = _zz_4654[15 : 0];
  assign _zz_359 = 1'b1;
  assign _zz_360 = 1'b1;
  assign _zz_1973 = ($signed(_zz_4671) - $signed(_zz_4672));
  assign _zz_361 = _zz_4673[15 : 0];
  assign _zz_1974 = ($signed(_zz_4674) + $signed(_zz_4675));
  assign _zz_362 = _zz_4676[15 : 0];
  assign _zz_363 = 1'b1;
  assign _zz_364 = 1'b1;
  assign _zz_1975 = ($signed(_zz_4693) - $signed(_zz_4694));
  assign _zz_365 = _zz_4695[15 : 0];
  assign _zz_1976 = ($signed(_zz_4696) + $signed(_zz_4697));
  assign _zz_366 = _zz_4698[15 : 0];
  assign _zz_367 = 1'b1;
  assign _zz_368 = 1'b1;
  assign _zz_1977 = ($signed(_zz_4715) - $signed(_zz_4716));
  assign _zz_369 = _zz_4717[15 : 0];
  assign _zz_1978 = ($signed(_zz_4718) + $signed(_zz_4719));
  assign _zz_370 = _zz_4720[15 : 0];
  assign _zz_371 = 1'b1;
  assign _zz_372 = 1'b1;
  assign _zz_1979 = ($signed(_zz_4737) - $signed(_zz_4738));
  assign _zz_373 = _zz_4739[15 : 0];
  assign _zz_1980 = ($signed(_zz_4740) + $signed(_zz_4741));
  assign _zz_374 = _zz_4742[15 : 0];
  assign _zz_375 = 1'b1;
  assign _zz_376 = 1'b1;
  assign _zz_1981 = ($signed(_zz_4759) - $signed(_zz_4760));
  assign _zz_377 = _zz_4761[15 : 0];
  assign _zz_1982 = ($signed(_zz_4762) + $signed(_zz_4763));
  assign _zz_378 = _zz_4764[15 : 0];
  assign _zz_379 = 1'b1;
  assign _zz_380 = 1'b1;
  assign _zz_1983 = ($signed(_zz_4781) - $signed(_zz_4782));
  assign _zz_381 = _zz_4783[15 : 0];
  assign _zz_1984 = ($signed(_zz_4784) + $signed(_zz_4785));
  assign _zz_382 = _zz_4786[15 : 0];
  assign _zz_383 = 1'b1;
  assign _zz_384 = 1'b1;
  assign _zz_1985 = ($signed(_zz_4803) - $signed(_zz_4804));
  assign _zz_385 = _zz_4805[15 : 0];
  assign _zz_1986 = ($signed(_zz_4806) + $signed(_zz_4807));
  assign _zz_386 = _zz_4808[15 : 0];
  assign _zz_387 = 1'b1;
  assign _zz_388 = 1'b1;
  assign _zz_1987 = ($signed(_zz_4825) - $signed(_zz_4826));
  assign _zz_389 = _zz_4827[15 : 0];
  assign _zz_1988 = ($signed(_zz_4828) + $signed(_zz_4829));
  assign _zz_390 = _zz_4830[15 : 0];
  assign _zz_391 = 1'b1;
  assign _zz_392 = 1'b1;
  assign _zz_1989 = ($signed(_zz_4847) - $signed(_zz_4848));
  assign _zz_393 = _zz_4849[15 : 0];
  assign _zz_1990 = ($signed(_zz_4850) + $signed(_zz_4851));
  assign _zz_394 = _zz_4852[15 : 0];
  assign _zz_395 = 1'b1;
  assign _zz_396 = 1'b1;
  assign _zz_1991 = ($signed(_zz_4869) - $signed(_zz_4870));
  assign _zz_397 = _zz_4871[15 : 0];
  assign _zz_1992 = ($signed(_zz_4872) + $signed(_zz_4873));
  assign _zz_398 = _zz_4874[15 : 0];
  assign _zz_399 = 1'b1;
  assign _zz_400 = 1'b1;
  assign _zz_1993 = ($signed(_zz_4891) - $signed(_zz_4892));
  assign _zz_401 = _zz_4893[15 : 0];
  assign _zz_1994 = ($signed(_zz_4894) + $signed(_zz_4895));
  assign _zz_402 = _zz_4896[15 : 0];
  assign _zz_403 = 1'b1;
  assign _zz_404 = 1'b1;
  assign _zz_1995 = ($signed(_zz_4913) - $signed(_zz_4914));
  assign _zz_405 = _zz_4915[15 : 0];
  assign _zz_1996 = ($signed(_zz_4916) + $signed(_zz_4917));
  assign _zz_406 = _zz_4918[15 : 0];
  assign _zz_407 = 1'b1;
  assign _zz_408 = 1'b1;
  assign _zz_1997 = ($signed(_zz_4935) - $signed(_zz_4936));
  assign _zz_409 = _zz_4937[15 : 0];
  assign _zz_1998 = ($signed(_zz_4938) + $signed(_zz_4939));
  assign _zz_410 = _zz_4940[15 : 0];
  assign _zz_411 = 1'b1;
  assign _zz_412 = 1'b1;
  assign _zz_1999 = ($signed(_zz_4957) - $signed(_zz_4958));
  assign _zz_413 = _zz_4959[15 : 0];
  assign _zz_2000 = ($signed(_zz_4960) + $signed(_zz_4961));
  assign _zz_414 = _zz_4962[15 : 0];
  assign _zz_415 = 1'b1;
  assign _zz_416 = 1'b1;
  assign _zz_2001 = ($signed(_zz_4979) - $signed(_zz_4980));
  assign _zz_417 = _zz_4981[15 : 0];
  assign _zz_2002 = ($signed(_zz_4982) + $signed(_zz_4983));
  assign _zz_418 = _zz_4984[15 : 0];
  assign _zz_419 = 1'b1;
  assign _zz_420 = 1'b1;
  assign _zz_2003 = ($signed(_zz_5001) - $signed(_zz_5002));
  assign _zz_421 = _zz_5003[15 : 0];
  assign _zz_2004 = ($signed(_zz_5004) + $signed(_zz_5005));
  assign _zz_422 = _zz_5006[15 : 0];
  assign _zz_423 = 1'b1;
  assign _zz_424 = 1'b1;
  assign _zz_2005 = ($signed(_zz_5023) - $signed(_zz_5024));
  assign _zz_425 = _zz_5025[15 : 0];
  assign _zz_2006 = ($signed(_zz_5026) + $signed(_zz_5027));
  assign _zz_426 = _zz_5028[15 : 0];
  assign _zz_427 = 1'b1;
  assign _zz_428 = 1'b1;
  assign _zz_2007 = ($signed(_zz_5045) - $signed(_zz_5046));
  assign _zz_429 = _zz_5047[15 : 0];
  assign _zz_2008 = ($signed(_zz_5048) + $signed(_zz_5049));
  assign _zz_430 = _zz_5050[15 : 0];
  assign _zz_431 = 1'b1;
  assign _zz_432 = 1'b1;
  assign _zz_2009 = ($signed(_zz_5067) - $signed(_zz_5068));
  assign _zz_433 = _zz_5069[15 : 0];
  assign _zz_2010 = ($signed(_zz_5070) + $signed(_zz_5071));
  assign _zz_434 = _zz_5072[15 : 0];
  assign _zz_435 = 1'b1;
  assign _zz_436 = 1'b1;
  assign _zz_2011 = ($signed(_zz_5089) - $signed(_zz_5090));
  assign _zz_437 = _zz_5091[15 : 0];
  assign _zz_2012 = ($signed(_zz_5092) + $signed(_zz_5093));
  assign _zz_438 = _zz_5094[15 : 0];
  assign _zz_439 = 1'b1;
  assign _zz_440 = 1'b1;
  assign _zz_2013 = ($signed(_zz_5111) - $signed(_zz_5112));
  assign _zz_441 = _zz_5113[15 : 0];
  assign _zz_2014 = ($signed(_zz_5114) + $signed(_zz_5115));
  assign _zz_442 = _zz_5116[15 : 0];
  assign _zz_443 = 1'b1;
  assign _zz_444 = 1'b1;
  assign _zz_2015 = ($signed(_zz_5133) - $signed(_zz_5134));
  assign _zz_445 = _zz_5135[15 : 0];
  assign _zz_2016 = ($signed(_zz_5136) + $signed(_zz_5137));
  assign _zz_446 = _zz_5138[15 : 0];
  assign _zz_447 = 1'b1;
  assign _zz_448 = 1'b1;
  assign _zz_2017 = ($signed(_zz_5155) - $signed(_zz_5156));
  assign _zz_449 = _zz_5157[15 : 0];
  assign _zz_2018 = ($signed(_zz_5158) + $signed(_zz_5159));
  assign _zz_450 = _zz_5160[15 : 0];
  assign _zz_451 = 1'b1;
  assign _zz_452 = 1'b1;
  assign _zz_2019 = ($signed(_zz_5177) - $signed(_zz_5178));
  assign _zz_453 = _zz_5179[15 : 0];
  assign _zz_2020 = ($signed(_zz_5180) + $signed(_zz_5181));
  assign _zz_454 = _zz_5182[15 : 0];
  assign _zz_455 = 1'b1;
  assign _zz_456 = 1'b1;
  assign _zz_2021 = ($signed(_zz_5199) - $signed(_zz_5200));
  assign _zz_457 = _zz_5201[15 : 0];
  assign _zz_2022 = ($signed(_zz_5202) + $signed(_zz_5203));
  assign _zz_458 = _zz_5204[15 : 0];
  assign _zz_459 = 1'b1;
  assign _zz_460 = 1'b1;
  assign _zz_2023 = ($signed(_zz_5221) - $signed(_zz_5222));
  assign _zz_461 = _zz_5223[15 : 0];
  assign _zz_2024 = ($signed(_zz_5224) + $signed(_zz_5225));
  assign _zz_462 = _zz_5226[15 : 0];
  assign _zz_463 = 1'b1;
  assign _zz_464 = 1'b1;
  assign _zz_2025 = ($signed(_zz_5243) - $signed(_zz_5244));
  assign _zz_465 = _zz_5245[15 : 0];
  assign _zz_2026 = ($signed(_zz_5246) + $signed(_zz_5247));
  assign _zz_466 = _zz_5248[15 : 0];
  assign _zz_467 = 1'b1;
  assign _zz_468 = 1'b1;
  assign _zz_2027 = ($signed(_zz_5265) - $signed(_zz_5266));
  assign _zz_469 = _zz_5267[15 : 0];
  assign _zz_2028 = ($signed(_zz_5268) + $signed(_zz_5269));
  assign _zz_470 = _zz_5270[15 : 0];
  assign _zz_471 = 1'b1;
  assign _zz_472 = 1'b1;
  assign _zz_2029 = ($signed(_zz_5287) - $signed(_zz_5288));
  assign _zz_473 = _zz_5289[15 : 0];
  assign _zz_2030 = ($signed(_zz_5290) + $signed(_zz_5291));
  assign _zz_474 = _zz_5292[15 : 0];
  assign _zz_475 = 1'b1;
  assign _zz_476 = 1'b1;
  assign _zz_2031 = ($signed(_zz_5309) - $signed(_zz_5310));
  assign _zz_477 = _zz_5311[15 : 0];
  assign _zz_2032 = ($signed(_zz_5312) + $signed(_zz_5313));
  assign _zz_478 = _zz_5314[15 : 0];
  assign _zz_479 = 1'b1;
  assign _zz_480 = 1'b1;
  assign _zz_2033 = ($signed(_zz_5331) - $signed(_zz_5332));
  assign _zz_481 = _zz_5333[15 : 0];
  assign _zz_2034 = ($signed(_zz_5334) + $signed(_zz_5335));
  assign _zz_482 = _zz_5336[15 : 0];
  assign _zz_483 = 1'b1;
  assign _zz_484 = 1'b1;
  assign _zz_2035 = ($signed(_zz_5353) - $signed(_zz_5354));
  assign _zz_485 = _zz_5355[15 : 0];
  assign _zz_2036 = ($signed(_zz_5356) + $signed(_zz_5357));
  assign _zz_486 = _zz_5358[15 : 0];
  assign _zz_487 = 1'b1;
  assign _zz_488 = 1'b1;
  assign _zz_2037 = ($signed(_zz_5375) - $signed(_zz_5376));
  assign _zz_489 = _zz_5377[15 : 0];
  assign _zz_2038 = ($signed(_zz_5378) + $signed(_zz_5379));
  assign _zz_490 = _zz_5380[15 : 0];
  assign _zz_491 = 1'b1;
  assign _zz_492 = 1'b1;
  assign _zz_2039 = ($signed(_zz_5397) - $signed(_zz_5398));
  assign _zz_493 = _zz_5399[15 : 0];
  assign _zz_2040 = ($signed(_zz_5400) + $signed(_zz_5401));
  assign _zz_494 = _zz_5402[15 : 0];
  assign _zz_495 = 1'b1;
  assign _zz_496 = 1'b1;
  assign _zz_2041 = ($signed(_zz_5419) - $signed(_zz_5420));
  assign _zz_497 = _zz_5421[15 : 0];
  assign _zz_2042 = ($signed(_zz_5422) + $signed(_zz_5423));
  assign _zz_498 = _zz_5424[15 : 0];
  assign _zz_499 = 1'b1;
  assign _zz_500 = 1'b1;
  assign _zz_2043 = ($signed(_zz_5441) - $signed(_zz_5442));
  assign _zz_501 = _zz_5443[15 : 0];
  assign _zz_2044 = ($signed(_zz_5444) + $signed(_zz_5445));
  assign _zz_502 = _zz_5446[15 : 0];
  assign _zz_503 = 1'b1;
  assign _zz_504 = 1'b1;
  assign _zz_2045 = ($signed(_zz_5463) - $signed(_zz_5464));
  assign _zz_505 = _zz_5465[15 : 0];
  assign _zz_2046 = ($signed(_zz_5466) + $signed(_zz_5467));
  assign _zz_506 = _zz_5468[15 : 0];
  assign _zz_507 = 1'b1;
  assign _zz_508 = 1'b1;
  assign _zz_2047 = ($signed(_zz_5485) - $signed(_zz_5486));
  assign _zz_509 = _zz_5487[15 : 0];
  assign _zz_2048 = ($signed(_zz_5488) + $signed(_zz_5489));
  assign _zz_510 = _zz_5490[15 : 0];
  assign _zz_511 = 1'b1;
  assign _zz_512 = 1'b1;
  assign _zz_2049 = ($signed(_zz_5507) - $signed(_zz_5508));
  assign _zz_513 = _zz_5509[15 : 0];
  assign _zz_2050 = ($signed(_zz_5510) + $signed(_zz_5511));
  assign _zz_514 = _zz_5512[15 : 0];
  assign _zz_515 = 1'b1;
  assign _zz_516 = 1'b1;
  assign _zz_2051 = ($signed(_zz_5529) - $signed(_zz_5530));
  assign _zz_517 = _zz_5531[15 : 0];
  assign _zz_2052 = ($signed(_zz_5532) + $signed(_zz_5533));
  assign _zz_518 = _zz_5534[15 : 0];
  assign _zz_519 = 1'b1;
  assign _zz_520 = 1'b1;
  assign _zz_2053 = ($signed(_zz_5551) - $signed(_zz_5552));
  assign _zz_521 = _zz_5553[15 : 0];
  assign _zz_2054 = ($signed(_zz_5554) + $signed(_zz_5555));
  assign _zz_522 = _zz_5556[15 : 0];
  assign _zz_523 = 1'b1;
  assign _zz_524 = 1'b1;
  assign _zz_2055 = ($signed(_zz_5573) - $signed(_zz_5574));
  assign _zz_525 = _zz_5575[15 : 0];
  assign _zz_2056 = ($signed(_zz_5576) + $signed(_zz_5577));
  assign _zz_526 = _zz_5578[15 : 0];
  assign _zz_527 = 1'b1;
  assign _zz_528 = 1'b1;
  assign _zz_2057 = ($signed(_zz_5595) - $signed(_zz_5596));
  assign _zz_529 = _zz_5597[15 : 0];
  assign _zz_2058 = ($signed(_zz_5598) + $signed(_zz_5599));
  assign _zz_530 = _zz_5600[15 : 0];
  assign _zz_531 = 1'b1;
  assign _zz_532 = 1'b1;
  assign _zz_2059 = ($signed(_zz_5617) - $signed(_zz_5618));
  assign _zz_533 = _zz_5619[15 : 0];
  assign _zz_2060 = ($signed(_zz_5620) + $signed(_zz_5621));
  assign _zz_534 = _zz_5622[15 : 0];
  assign _zz_535 = 1'b1;
  assign _zz_536 = 1'b1;
  assign _zz_2061 = ($signed(_zz_5639) - $signed(_zz_5640));
  assign _zz_537 = _zz_5641[15 : 0];
  assign _zz_2062 = ($signed(_zz_5642) + $signed(_zz_5643));
  assign _zz_538 = _zz_5644[15 : 0];
  assign _zz_539 = 1'b1;
  assign _zz_540 = 1'b1;
  assign _zz_2063 = ($signed(_zz_5661) - $signed(_zz_5662));
  assign _zz_541 = _zz_5663[15 : 0];
  assign _zz_2064 = ($signed(_zz_5664) + $signed(_zz_5665));
  assign _zz_542 = _zz_5666[15 : 0];
  assign _zz_543 = 1'b1;
  assign _zz_544 = 1'b1;
  assign _zz_2065 = ($signed(_zz_5683) - $signed(_zz_5684));
  assign _zz_545 = _zz_5685[15 : 0];
  assign _zz_2066 = ($signed(_zz_5686) + $signed(_zz_5687));
  assign _zz_546 = _zz_5688[15 : 0];
  assign _zz_547 = 1'b1;
  assign _zz_548 = 1'b1;
  assign _zz_2067 = ($signed(_zz_5705) - $signed(_zz_5706));
  assign _zz_549 = _zz_5707[15 : 0];
  assign _zz_2068 = ($signed(_zz_5708) + $signed(_zz_5709));
  assign _zz_550 = _zz_5710[15 : 0];
  assign _zz_551 = 1'b1;
  assign _zz_552 = 1'b1;
  assign _zz_2069 = ($signed(_zz_5727) - $signed(_zz_5728));
  assign _zz_553 = _zz_5729[15 : 0];
  assign _zz_2070 = ($signed(_zz_5730) + $signed(_zz_5731));
  assign _zz_554 = _zz_5732[15 : 0];
  assign _zz_555 = 1'b1;
  assign _zz_556 = 1'b1;
  assign _zz_2071 = ($signed(_zz_5749) - $signed(_zz_5750));
  assign _zz_557 = _zz_5751[15 : 0];
  assign _zz_2072 = ($signed(_zz_5752) + $signed(_zz_5753));
  assign _zz_558 = _zz_5754[15 : 0];
  assign _zz_559 = 1'b1;
  assign _zz_560 = 1'b1;
  assign _zz_2073 = ($signed(_zz_5771) - $signed(_zz_5772));
  assign _zz_561 = _zz_5773[15 : 0];
  assign _zz_2074 = ($signed(_zz_5774) + $signed(_zz_5775));
  assign _zz_562 = _zz_5776[15 : 0];
  assign _zz_563 = 1'b1;
  assign _zz_564 = 1'b1;
  assign _zz_2075 = ($signed(_zz_5793) - $signed(_zz_5794));
  assign _zz_565 = _zz_5795[15 : 0];
  assign _zz_2076 = ($signed(_zz_5796) + $signed(_zz_5797));
  assign _zz_566 = _zz_5798[15 : 0];
  assign _zz_567 = 1'b1;
  assign _zz_568 = 1'b1;
  assign _zz_2077 = ($signed(_zz_5815) - $signed(_zz_5816));
  assign _zz_569 = _zz_5817[15 : 0];
  assign _zz_2078 = ($signed(_zz_5818) + $signed(_zz_5819));
  assign _zz_570 = _zz_5820[15 : 0];
  assign _zz_571 = 1'b1;
  assign _zz_572 = 1'b1;
  assign _zz_2079 = ($signed(_zz_5837) - $signed(_zz_5838));
  assign _zz_573 = _zz_5839[15 : 0];
  assign _zz_2080 = ($signed(_zz_5840) + $signed(_zz_5841));
  assign _zz_574 = _zz_5842[15 : 0];
  assign _zz_575 = 1'b1;
  assign _zz_576 = 1'b1;
  assign _zz_2081 = ($signed(_zz_5859) - $signed(_zz_5860));
  assign _zz_577 = _zz_5861[15 : 0];
  assign _zz_2082 = ($signed(_zz_5862) + $signed(_zz_5863));
  assign _zz_578 = _zz_5864[15 : 0];
  assign _zz_579 = 1'b1;
  assign _zz_580 = 1'b1;
  assign _zz_2083 = ($signed(_zz_5881) - $signed(_zz_5882));
  assign _zz_581 = _zz_5883[15 : 0];
  assign _zz_2084 = ($signed(_zz_5884) + $signed(_zz_5885));
  assign _zz_582 = _zz_5886[15 : 0];
  assign _zz_583 = 1'b1;
  assign _zz_584 = 1'b1;
  assign _zz_2085 = ($signed(_zz_5903) - $signed(_zz_5904));
  assign _zz_585 = _zz_5905[15 : 0];
  assign _zz_2086 = ($signed(_zz_5906) + $signed(_zz_5907));
  assign _zz_586 = _zz_5908[15 : 0];
  assign _zz_587 = 1'b1;
  assign _zz_588 = 1'b1;
  assign _zz_2087 = ($signed(_zz_5925) - $signed(_zz_5926));
  assign _zz_589 = _zz_5927[15 : 0];
  assign _zz_2088 = ($signed(_zz_5928) + $signed(_zz_5929));
  assign _zz_590 = _zz_5930[15 : 0];
  assign _zz_591 = 1'b1;
  assign _zz_592 = 1'b1;
  assign _zz_2089 = ($signed(_zz_5947) - $signed(_zz_5948));
  assign _zz_593 = _zz_5949[15 : 0];
  assign _zz_2090 = ($signed(_zz_5950) + $signed(_zz_5951));
  assign _zz_594 = _zz_5952[15 : 0];
  assign _zz_595 = 1'b1;
  assign _zz_596 = 1'b1;
  assign _zz_2091 = ($signed(_zz_5969) - $signed(_zz_5970));
  assign _zz_597 = _zz_5971[15 : 0];
  assign _zz_2092 = ($signed(_zz_5972) + $signed(_zz_5973));
  assign _zz_598 = _zz_5974[15 : 0];
  assign _zz_599 = 1'b1;
  assign _zz_600 = 1'b1;
  assign _zz_2093 = ($signed(_zz_5991) - $signed(_zz_5992));
  assign _zz_601 = _zz_5993[15 : 0];
  assign _zz_2094 = ($signed(_zz_5994) + $signed(_zz_5995));
  assign _zz_602 = _zz_5996[15 : 0];
  assign _zz_603 = 1'b1;
  assign _zz_604 = 1'b1;
  assign _zz_2095 = ($signed(_zz_6013) - $signed(_zz_6014));
  assign _zz_605 = _zz_6015[15 : 0];
  assign _zz_2096 = ($signed(_zz_6016) + $signed(_zz_6017));
  assign _zz_606 = _zz_6018[15 : 0];
  assign _zz_607 = 1'b1;
  assign _zz_608 = 1'b1;
  assign _zz_2097 = ($signed(_zz_6035) - $signed(_zz_6036));
  assign _zz_609 = _zz_6037[15 : 0];
  assign _zz_2098 = ($signed(_zz_6038) + $signed(_zz_6039));
  assign _zz_610 = _zz_6040[15 : 0];
  assign _zz_611 = 1'b1;
  assign _zz_612 = 1'b1;
  assign _zz_2099 = ($signed(_zz_6057) - $signed(_zz_6058));
  assign _zz_613 = _zz_6059[15 : 0];
  assign _zz_2100 = ($signed(_zz_6060) + $signed(_zz_6061));
  assign _zz_614 = _zz_6062[15 : 0];
  assign _zz_615 = 1'b1;
  assign _zz_616 = 1'b1;
  assign _zz_2101 = ($signed(_zz_6079) - $signed(_zz_6080));
  assign _zz_617 = _zz_6081[15 : 0];
  assign _zz_2102 = ($signed(_zz_6082) + $signed(_zz_6083));
  assign _zz_618 = _zz_6084[15 : 0];
  assign _zz_619 = 1'b1;
  assign _zz_620 = 1'b1;
  assign _zz_2103 = ($signed(_zz_6101) - $signed(_zz_6102));
  assign _zz_621 = _zz_6103[15 : 0];
  assign _zz_2104 = ($signed(_zz_6104) + $signed(_zz_6105));
  assign _zz_622 = _zz_6106[15 : 0];
  assign _zz_623 = 1'b1;
  assign _zz_624 = 1'b1;
  assign _zz_2105 = ($signed(_zz_6123) - $signed(_zz_6124));
  assign _zz_625 = _zz_6125[15 : 0];
  assign _zz_2106 = ($signed(_zz_6126) + $signed(_zz_6127));
  assign _zz_626 = _zz_6128[15 : 0];
  assign _zz_627 = 1'b1;
  assign _zz_628 = 1'b1;
  assign _zz_2107 = ($signed(_zz_6145) - $signed(_zz_6146));
  assign _zz_629 = _zz_6147[15 : 0];
  assign _zz_2108 = ($signed(_zz_6148) + $signed(_zz_6149));
  assign _zz_630 = _zz_6150[15 : 0];
  assign _zz_631 = 1'b1;
  assign _zz_632 = 1'b1;
  assign _zz_2109 = ($signed(_zz_6167) - $signed(_zz_6168));
  assign _zz_633 = _zz_6169[15 : 0];
  assign _zz_2110 = ($signed(_zz_6170) + $signed(_zz_6171));
  assign _zz_634 = _zz_6172[15 : 0];
  assign _zz_635 = 1'b1;
  assign _zz_636 = 1'b1;
  assign _zz_2111 = ($signed(_zz_6189) - $signed(_zz_6190));
  assign _zz_637 = _zz_6191[15 : 0];
  assign _zz_2112 = ($signed(_zz_6192) + $signed(_zz_6193));
  assign _zz_638 = _zz_6194[15 : 0];
  assign _zz_639 = 1'b1;
  assign _zz_640 = 1'b1;
  assign _zz_2113 = ($signed(_zz_6211) - $signed(_zz_6212));
  assign _zz_641 = _zz_6213[15 : 0];
  assign _zz_2114 = ($signed(_zz_6214) + $signed(_zz_6215));
  assign _zz_642 = _zz_6216[15 : 0];
  assign _zz_643 = 1'b1;
  assign _zz_644 = 1'b1;
  assign _zz_2115 = ($signed(_zz_6233) - $signed(_zz_6234));
  assign _zz_645 = _zz_6235[15 : 0];
  assign _zz_2116 = ($signed(_zz_6236) + $signed(_zz_6237));
  assign _zz_646 = _zz_6238[15 : 0];
  assign _zz_647 = 1'b1;
  assign _zz_648 = 1'b1;
  assign _zz_2117 = ($signed(_zz_6255) - $signed(_zz_6256));
  assign _zz_649 = _zz_6257[15 : 0];
  assign _zz_2118 = ($signed(_zz_6258) + $signed(_zz_6259));
  assign _zz_650 = _zz_6260[15 : 0];
  assign _zz_651 = 1'b1;
  assign _zz_652 = 1'b1;
  assign _zz_2119 = ($signed(_zz_6277) - $signed(_zz_6278));
  assign _zz_653 = _zz_6279[15 : 0];
  assign _zz_2120 = ($signed(_zz_6280) + $signed(_zz_6281));
  assign _zz_654 = _zz_6282[15 : 0];
  assign _zz_655 = 1'b1;
  assign _zz_656 = 1'b1;
  assign _zz_2121 = ($signed(_zz_6299) - $signed(_zz_6300));
  assign _zz_657 = _zz_6301[15 : 0];
  assign _zz_2122 = ($signed(_zz_6302) + $signed(_zz_6303));
  assign _zz_658 = _zz_6304[15 : 0];
  assign _zz_659 = 1'b1;
  assign _zz_660 = 1'b1;
  assign _zz_2123 = ($signed(_zz_6321) - $signed(_zz_6322));
  assign _zz_661 = _zz_6323[15 : 0];
  assign _zz_2124 = ($signed(_zz_6324) + $signed(_zz_6325));
  assign _zz_662 = _zz_6326[15 : 0];
  assign _zz_663 = 1'b1;
  assign _zz_664 = 1'b1;
  assign _zz_2125 = ($signed(_zz_6343) - $signed(_zz_6344));
  assign _zz_665 = _zz_6345[15 : 0];
  assign _zz_2126 = ($signed(_zz_6346) + $signed(_zz_6347));
  assign _zz_666 = _zz_6348[15 : 0];
  assign _zz_667 = 1'b1;
  assign _zz_668 = 1'b1;
  assign _zz_2127 = ($signed(_zz_6365) - $signed(_zz_6366));
  assign _zz_669 = _zz_6367[15 : 0];
  assign _zz_2128 = ($signed(_zz_6368) + $signed(_zz_6369));
  assign _zz_670 = _zz_6370[15 : 0];
  assign _zz_671 = 1'b1;
  assign _zz_672 = 1'b1;
  assign _zz_2129 = ($signed(_zz_6387) - $signed(_zz_6388));
  assign _zz_673 = _zz_6389[15 : 0];
  assign _zz_2130 = ($signed(_zz_6390) + $signed(_zz_6391));
  assign _zz_674 = _zz_6392[15 : 0];
  assign _zz_675 = 1'b1;
  assign _zz_676 = 1'b1;
  assign _zz_2131 = ($signed(_zz_6409) - $signed(_zz_6410));
  assign _zz_677 = _zz_6411[15 : 0];
  assign _zz_2132 = ($signed(_zz_6412) + $signed(_zz_6413));
  assign _zz_678 = _zz_6414[15 : 0];
  assign _zz_679 = 1'b1;
  assign _zz_680 = 1'b1;
  assign _zz_2133 = ($signed(_zz_6431) - $signed(_zz_6432));
  assign _zz_681 = _zz_6433[15 : 0];
  assign _zz_2134 = ($signed(_zz_6434) + $signed(_zz_6435));
  assign _zz_682 = _zz_6436[15 : 0];
  assign _zz_683 = 1'b1;
  assign _zz_684 = 1'b1;
  assign _zz_2135 = ($signed(_zz_6453) - $signed(_zz_6454));
  assign _zz_685 = _zz_6455[15 : 0];
  assign _zz_2136 = ($signed(_zz_6456) + $signed(_zz_6457));
  assign _zz_686 = _zz_6458[15 : 0];
  assign _zz_687 = 1'b1;
  assign _zz_688 = 1'b1;
  assign _zz_2137 = ($signed(_zz_6475) - $signed(_zz_6476));
  assign _zz_689 = _zz_6477[15 : 0];
  assign _zz_2138 = ($signed(_zz_6478) + $signed(_zz_6479));
  assign _zz_690 = _zz_6480[15 : 0];
  assign _zz_691 = 1'b1;
  assign _zz_692 = 1'b1;
  assign _zz_2139 = ($signed(_zz_6497) - $signed(_zz_6498));
  assign _zz_693 = _zz_6499[15 : 0];
  assign _zz_2140 = ($signed(_zz_6500) + $signed(_zz_6501));
  assign _zz_694 = _zz_6502[15 : 0];
  assign _zz_695 = 1'b1;
  assign _zz_696 = 1'b1;
  assign _zz_2141 = ($signed(_zz_6519) - $signed(_zz_6520));
  assign _zz_697 = _zz_6521[15 : 0];
  assign _zz_2142 = ($signed(_zz_6522) + $signed(_zz_6523));
  assign _zz_698 = _zz_6524[15 : 0];
  assign _zz_699 = 1'b1;
  assign _zz_700 = 1'b1;
  assign _zz_2143 = ($signed(_zz_6541) - $signed(_zz_6542));
  assign _zz_701 = _zz_6543[15 : 0];
  assign _zz_2144 = ($signed(_zz_6544) + $signed(_zz_6545));
  assign _zz_702 = _zz_6546[15 : 0];
  assign _zz_703 = 1'b1;
  assign _zz_704 = 1'b1;
  assign _zz_2145 = ($signed(_zz_6563) - $signed(_zz_6564));
  assign _zz_705 = _zz_6565[15 : 0];
  assign _zz_2146 = ($signed(_zz_6566) + $signed(_zz_6567));
  assign _zz_706 = _zz_6568[15 : 0];
  assign _zz_707 = 1'b1;
  assign _zz_708 = 1'b1;
  assign _zz_2147 = ($signed(_zz_6585) - $signed(_zz_6586));
  assign _zz_709 = _zz_6587[15 : 0];
  assign _zz_2148 = ($signed(_zz_6588) + $signed(_zz_6589));
  assign _zz_710 = _zz_6590[15 : 0];
  assign _zz_711 = 1'b1;
  assign _zz_712 = 1'b1;
  assign _zz_2149 = ($signed(_zz_6607) - $signed(_zz_6608));
  assign _zz_713 = _zz_6609[15 : 0];
  assign _zz_2150 = ($signed(_zz_6610) + $signed(_zz_6611));
  assign _zz_714 = _zz_6612[15 : 0];
  assign _zz_715 = 1'b1;
  assign _zz_716 = 1'b1;
  assign _zz_2151 = ($signed(_zz_6629) - $signed(_zz_6630));
  assign _zz_717 = _zz_6631[15 : 0];
  assign _zz_2152 = ($signed(_zz_6632) + $signed(_zz_6633));
  assign _zz_718 = _zz_6634[15 : 0];
  assign _zz_719 = 1'b1;
  assign _zz_720 = 1'b1;
  assign _zz_2153 = ($signed(_zz_6651) - $signed(_zz_6652));
  assign _zz_721 = _zz_6653[15 : 0];
  assign _zz_2154 = ($signed(_zz_6654) + $signed(_zz_6655));
  assign _zz_722 = _zz_6656[15 : 0];
  assign _zz_723 = 1'b1;
  assign _zz_724 = 1'b1;
  assign _zz_2155 = ($signed(_zz_6673) - $signed(_zz_6674));
  assign _zz_725 = _zz_6675[15 : 0];
  assign _zz_2156 = ($signed(_zz_6676) + $signed(_zz_6677));
  assign _zz_726 = _zz_6678[15 : 0];
  assign _zz_727 = 1'b1;
  assign _zz_728 = 1'b1;
  assign _zz_2157 = ($signed(_zz_6695) - $signed(_zz_6696));
  assign _zz_729 = _zz_6697[15 : 0];
  assign _zz_2158 = ($signed(_zz_6698) + $signed(_zz_6699));
  assign _zz_730 = _zz_6700[15 : 0];
  assign _zz_731 = 1'b1;
  assign _zz_732 = 1'b1;
  assign _zz_2159 = ($signed(_zz_6717) - $signed(_zz_6718));
  assign _zz_733 = _zz_6719[15 : 0];
  assign _zz_2160 = ($signed(_zz_6720) + $signed(_zz_6721));
  assign _zz_734 = _zz_6722[15 : 0];
  assign _zz_735 = 1'b1;
  assign _zz_736 = 1'b1;
  assign _zz_2161 = ($signed(_zz_6739) - $signed(_zz_6740));
  assign _zz_737 = _zz_6741[15 : 0];
  assign _zz_2162 = ($signed(_zz_6742) + $signed(_zz_6743));
  assign _zz_738 = _zz_6744[15 : 0];
  assign _zz_739 = 1'b1;
  assign _zz_740 = 1'b1;
  assign _zz_2163 = ($signed(_zz_6761) - $signed(_zz_6762));
  assign _zz_741 = _zz_6763[15 : 0];
  assign _zz_2164 = ($signed(_zz_6764) + $signed(_zz_6765));
  assign _zz_742 = _zz_6766[15 : 0];
  assign _zz_743 = 1'b1;
  assign _zz_744 = 1'b1;
  assign _zz_2165 = ($signed(_zz_6783) - $signed(_zz_6784));
  assign _zz_745 = _zz_6785[15 : 0];
  assign _zz_2166 = ($signed(_zz_6786) + $signed(_zz_6787));
  assign _zz_746 = _zz_6788[15 : 0];
  assign _zz_747 = 1'b1;
  assign _zz_748 = 1'b1;
  assign _zz_2167 = ($signed(_zz_6805) - $signed(_zz_6806));
  assign _zz_749 = _zz_6807[15 : 0];
  assign _zz_2168 = ($signed(_zz_6808) + $signed(_zz_6809));
  assign _zz_750 = _zz_6810[15 : 0];
  assign _zz_751 = 1'b1;
  assign _zz_752 = 1'b1;
  assign _zz_2169 = ($signed(_zz_6827) - $signed(_zz_6828));
  assign _zz_753 = _zz_6829[15 : 0];
  assign _zz_2170 = ($signed(_zz_6830) + $signed(_zz_6831));
  assign _zz_754 = _zz_6832[15 : 0];
  assign _zz_755 = 1'b1;
  assign _zz_756 = 1'b1;
  assign _zz_2171 = ($signed(_zz_6849) - $signed(_zz_6850));
  assign _zz_757 = _zz_6851[15 : 0];
  assign _zz_2172 = ($signed(_zz_6852) + $signed(_zz_6853));
  assign _zz_758 = _zz_6854[15 : 0];
  assign _zz_759 = 1'b1;
  assign _zz_760 = 1'b1;
  assign _zz_2173 = ($signed(_zz_6871) - $signed(_zz_6872));
  assign _zz_761 = _zz_6873[15 : 0];
  assign _zz_2174 = ($signed(_zz_6874) + $signed(_zz_6875));
  assign _zz_762 = _zz_6876[15 : 0];
  assign _zz_763 = 1'b1;
  assign _zz_764 = 1'b1;
  assign _zz_2175 = ($signed(_zz_6893) - $signed(_zz_6894));
  assign _zz_765 = _zz_6895[15 : 0];
  assign _zz_2176 = ($signed(_zz_6896) + $signed(_zz_6897));
  assign _zz_766 = _zz_6898[15 : 0];
  assign _zz_767 = 1'b1;
  assign _zz_768 = 1'b1;
  assign _zz_2177 = ($signed(_zz_6915) - $signed(_zz_6916));
  assign _zz_769 = _zz_6917[15 : 0];
  assign _zz_2178 = ($signed(_zz_6918) + $signed(_zz_6919));
  assign _zz_770 = _zz_6920[15 : 0];
  assign _zz_771 = 1'b1;
  assign _zz_772 = 1'b1;
  assign _zz_2179 = ($signed(_zz_6937) - $signed(_zz_6938));
  assign _zz_773 = _zz_6939[15 : 0];
  assign _zz_2180 = ($signed(_zz_6940) + $signed(_zz_6941));
  assign _zz_774 = _zz_6942[15 : 0];
  assign _zz_775 = 1'b1;
  assign _zz_776 = 1'b1;
  assign _zz_2181 = ($signed(_zz_6959) - $signed(_zz_6960));
  assign _zz_777 = _zz_6961[15 : 0];
  assign _zz_2182 = ($signed(_zz_6962) + $signed(_zz_6963));
  assign _zz_778 = _zz_6964[15 : 0];
  assign _zz_779 = 1'b1;
  assign _zz_780 = 1'b1;
  assign _zz_2183 = ($signed(_zz_6981) - $signed(_zz_6982));
  assign _zz_781 = _zz_6983[15 : 0];
  assign _zz_2184 = ($signed(_zz_6984) + $signed(_zz_6985));
  assign _zz_782 = _zz_6986[15 : 0];
  assign _zz_783 = 1'b1;
  assign _zz_784 = 1'b1;
  assign _zz_2185 = ($signed(_zz_7003) - $signed(_zz_7004));
  assign _zz_785 = _zz_7005[15 : 0];
  assign _zz_2186 = ($signed(_zz_7006) + $signed(_zz_7007));
  assign _zz_786 = _zz_7008[15 : 0];
  assign _zz_787 = 1'b1;
  assign _zz_788 = 1'b1;
  assign _zz_2187 = ($signed(_zz_7025) - $signed(_zz_7026));
  assign _zz_789 = _zz_7027[15 : 0];
  assign _zz_2188 = ($signed(_zz_7028) + $signed(_zz_7029));
  assign _zz_790 = _zz_7030[15 : 0];
  assign _zz_791 = 1'b1;
  assign _zz_792 = 1'b1;
  assign _zz_2189 = ($signed(_zz_7047) - $signed(_zz_7048));
  assign _zz_793 = _zz_7049[15 : 0];
  assign _zz_2190 = ($signed(_zz_7050) + $signed(_zz_7051));
  assign _zz_794 = _zz_7052[15 : 0];
  assign _zz_795 = 1'b1;
  assign _zz_796 = 1'b1;
  assign _zz_2191 = ($signed(_zz_7069) - $signed(_zz_7070));
  assign _zz_797 = _zz_7071[15 : 0];
  assign _zz_2192 = ($signed(_zz_7072) + $signed(_zz_7073));
  assign _zz_798 = _zz_7074[15 : 0];
  assign _zz_799 = 1'b1;
  assign _zz_800 = 1'b1;
  assign _zz_2193 = ($signed(_zz_7091) - $signed(_zz_7092));
  assign _zz_801 = _zz_7093[15 : 0];
  assign _zz_2194 = ($signed(_zz_7094) + $signed(_zz_7095));
  assign _zz_802 = _zz_7096[15 : 0];
  assign _zz_803 = 1'b1;
  assign _zz_804 = 1'b1;
  assign _zz_2195 = ($signed(_zz_7113) - $signed(_zz_7114));
  assign _zz_805 = _zz_7115[15 : 0];
  assign _zz_2196 = ($signed(_zz_7116) + $signed(_zz_7117));
  assign _zz_806 = _zz_7118[15 : 0];
  assign _zz_807 = 1'b1;
  assign _zz_808 = 1'b1;
  assign _zz_2197 = ($signed(_zz_7135) - $signed(_zz_7136));
  assign _zz_809 = _zz_7137[15 : 0];
  assign _zz_2198 = ($signed(_zz_7138) + $signed(_zz_7139));
  assign _zz_810 = _zz_7140[15 : 0];
  assign _zz_811 = 1'b1;
  assign _zz_812 = 1'b1;
  assign _zz_2199 = ($signed(_zz_7157) - $signed(_zz_7158));
  assign _zz_813 = _zz_7159[15 : 0];
  assign _zz_2200 = ($signed(_zz_7160) + $signed(_zz_7161));
  assign _zz_814 = _zz_7162[15 : 0];
  assign _zz_815 = 1'b1;
  assign _zz_816 = 1'b1;
  assign _zz_2201 = ($signed(_zz_7179) - $signed(_zz_7180));
  assign _zz_817 = _zz_7181[15 : 0];
  assign _zz_2202 = ($signed(_zz_7182) + $signed(_zz_7183));
  assign _zz_818 = _zz_7184[15 : 0];
  assign _zz_819 = 1'b1;
  assign _zz_820 = 1'b1;
  assign _zz_2203 = ($signed(_zz_7201) - $signed(_zz_7202));
  assign _zz_821 = _zz_7203[15 : 0];
  assign _zz_2204 = ($signed(_zz_7204) + $signed(_zz_7205));
  assign _zz_822 = _zz_7206[15 : 0];
  assign _zz_823 = 1'b1;
  assign _zz_824 = 1'b1;
  assign _zz_2205 = ($signed(_zz_7223) - $signed(_zz_7224));
  assign _zz_825 = _zz_7225[15 : 0];
  assign _zz_2206 = ($signed(_zz_7226) + $signed(_zz_7227));
  assign _zz_826 = _zz_7228[15 : 0];
  assign _zz_827 = 1'b1;
  assign _zz_828 = 1'b1;
  assign _zz_2207 = ($signed(_zz_7245) - $signed(_zz_7246));
  assign _zz_829 = _zz_7247[15 : 0];
  assign _zz_2208 = ($signed(_zz_7248) + $signed(_zz_7249));
  assign _zz_830 = _zz_7250[15 : 0];
  assign _zz_831 = 1'b1;
  assign _zz_832 = 1'b1;
  assign _zz_2209 = ($signed(_zz_7267) - $signed(_zz_7268));
  assign _zz_833 = _zz_7269[15 : 0];
  assign _zz_2210 = ($signed(_zz_7270) + $signed(_zz_7271));
  assign _zz_834 = _zz_7272[15 : 0];
  assign _zz_835 = 1'b1;
  assign _zz_836 = 1'b1;
  assign _zz_2211 = ($signed(_zz_7289) - $signed(_zz_7290));
  assign _zz_837 = _zz_7291[15 : 0];
  assign _zz_2212 = ($signed(_zz_7292) + $signed(_zz_7293));
  assign _zz_838 = _zz_7294[15 : 0];
  assign _zz_839 = 1'b1;
  assign _zz_840 = 1'b1;
  assign _zz_2213 = ($signed(_zz_7311) - $signed(_zz_7312));
  assign _zz_841 = _zz_7313[15 : 0];
  assign _zz_2214 = ($signed(_zz_7314) + $signed(_zz_7315));
  assign _zz_842 = _zz_7316[15 : 0];
  assign _zz_843 = 1'b1;
  assign _zz_844 = 1'b1;
  assign _zz_2215 = ($signed(_zz_7333) - $signed(_zz_7334));
  assign _zz_845 = _zz_7335[15 : 0];
  assign _zz_2216 = ($signed(_zz_7336) + $signed(_zz_7337));
  assign _zz_846 = _zz_7338[15 : 0];
  assign _zz_847 = 1'b1;
  assign _zz_848 = 1'b1;
  assign _zz_2217 = ($signed(_zz_7355) - $signed(_zz_7356));
  assign _zz_849 = _zz_7357[15 : 0];
  assign _zz_2218 = ($signed(_zz_7358) + $signed(_zz_7359));
  assign _zz_850 = _zz_7360[15 : 0];
  assign _zz_851 = 1'b1;
  assign _zz_852 = 1'b1;
  assign _zz_2219 = ($signed(_zz_7377) - $signed(_zz_7378));
  assign _zz_853 = _zz_7379[15 : 0];
  assign _zz_2220 = ($signed(_zz_7380) + $signed(_zz_7381));
  assign _zz_854 = _zz_7382[15 : 0];
  assign _zz_855 = 1'b1;
  assign _zz_856 = 1'b1;
  assign _zz_2221 = ($signed(_zz_7399) - $signed(_zz_7400));
  assign _zz_857 = _zz_7401[15 : 0];
  assign _zz_2222 = ($signed(_zz_7402) + $signed(_zz_7403));
  assign _zz_858 = _zz_7404[15 : 0];
  assign _zz_859 = 1'b1;
  assign _zz_860 = 1'b1;
  assign _zz_2223 = ($signed(_zz_7421) - $signed(_zz_7422));
  assign _zz_861 = _zz_7423[15 : 0];
  assign _zz_2224 = ($signed(_zz_7424) + $signed(_zz_7425));
  assign _zz_862 = _zz_7426[15 : 0];
  assign _zz_863 = 1'b1;
  assign _zz_864 = 1'b1;
  assign _zz_2225 = ($signed(_zz_7443) - $signed(_zz_7444));
  assign _zz_865 = _zz_7445[15 : 0];
  assign _zz_2226 = ($signed(_zz_7446) + $signed(_zz_7447));
  assign _zz_866 = _zz_7448[15 : 0];
  assign _zz_867 = 1'b1;
  assign _zz_868 = 1'b1;
  assign _zz_2227 = ($signed(_zz_7465) - $signed(_zz_7466));
  assign _zz_869 = _zz_7467[15 : 0];
  assign _zz_2228 = ($signed(_zz_7468) + $signed(_zz_7469));
  assign _zz_870 = _zz_7470[15 : 0];
  assign _zz_871 = 1'b1;
  assign _zz_872 = 1'b1;
  assign _zz_2229 = ($signed(_zz_7487) - $signed(_zz_7488));
  assign _zz_873 = _zz_7489[15 : 0];
  assign _zz_2230 = ($signed(_zz_7490) + $signed(_zz_7491));
  assign _zz_874 = _zz_7492[15 : 0];
  assign _zz_875 = 1'b1;
  assign _zz_876 = 1'b1;
  assign _zz_2231 = ($signed(_zz_7509) - $signed(_zz_7510));
  assign _zz_877 = _zz_7511[15 : 0];
  assign _zz_2232 = ($signed(_zz_7512) + $signed(_zz_7513));
  assign _zz_878 = _zz_7514[15 : 0];
  assign _zz_879 = 1'b1;
  assign _zz_880 = 1'b1;
  assign _zz_2233 = ($signed(_zz_7531) - $signed(_zz_7532));
  assign _zz_881 = _zz_7533[15 : 0];
  assign _zz_2234 = ($signed(_zz_7534) + $signed(_zz_7535));
  assign _zz_882 = _zz_7536[15 : 0];
  assign _zz_883 = 1'b1;
  assign _zz_884 = 1'b1;
  assign _zz_2235 = ($signed(_zz_7553) - $signed(_zz_7554));
  assign _zz_885 = _zz_7555[15 : 0];
  assign _zz_2236 = ($signed(_zz_7556) + $signed(_zz_7557));
  assign _zz_886 = _zz_7558[15 : 0];
  assign _zz_887 = 1'b1;
  assign _zz_888 = 1'b1;
  assign _zz_2237 = ($signed(_zz_7575) - $signed(_zz_7576));
  assign _zz_889 = _zz_7577[15 : 0];
  assign _zz_2238 = ($signed(_zz_7578) + $signed(_zz_7579));
  assign _zz_890 = _zz_7580[15 : 0];
  assign _zz_891 = 1'b1;
  assign _zz_892 = 1'b1;
  assign _zz_2239 = ($signed(_zz_7597) - $signed(_zz_7598));
  assign _zz_893 = _zz_7599[15 : 0];
  assign _zz_2240 = ($signed(_zz_7600) + $signed(_zz_7601));
  assign _zz_894 = _zz_7602[15 : 0];
  assign _zz_895 = 1'b1;
  assign _zz_896 = 1'b1;
  assign _zz_2241 = ($signed(_zz_7619) - $signed(_zz_7620));
  assign _zz_897 = _zz_7621[15 : 0];
  assign _zz_2242 = ($signed(_zz_7622) + $signed(_zz_7623));
  assign _zz_898 = _zz_7624[15 : 0];
  assign _zz_899 = 1'b1;
  assign _zz_900 = 1'b1;
  assign _zz_2243 = ($signed(_zz_7641) - $signed(_zz_7642));
  assign _zz_901 = _zz_7643[15 : 0];
  assign _zz_2244 = ($signed(_zz_7644) + $signed(_zz_7645));
  assign _zz_902 = _zz_7646[15 : 0];
  assign _zz_903 = 1'b1;
  assign _zz_904 = 1'b1;
  assign _zz_2245 = ($signed(_zz_7663) - $signed(_zz_7664));
  assign _zz_905 = _zz_7665[15 : 0];
  assign _zz_2246 = ($signed(_zz_7666) + $signed(_zz_7667));
  assign _zz_906 = _zz_7668[15 : 0];
  assign _zz_907 = 1'b1;
  assign _zz_908 = 1'b1;
  assign _zz_2247 = ($signed(_zz_7685) - $signed(_zz_7686));
  assign _zz_909 = _zz_7687[15 : 0];
  assign _zz_2248 = ($signed(_zz_7688) + $signed(_zz_7689));
  assign _zz_910 = _zz_7690[15 : 0];
  assign _zz_911 = 1'b1;
  assign _zz_912 = 1'b1;
  assign _zz_2249 = ($signed(_zz_7707) - $signed(_zz_7708));
  assign _zz_913 = _zz_7709[15 : 0];
  assign _zz_2250 = ($signed(_zz_7710) + $signed(_zz_7711));
  assign _zz_914 = _zz_7712[15 : 0];
  assign _zz_915 = 1'b1;
  assign _zz_916 = 1'b1;
  assign _zz_2251 = ($signed(_zz_7729) - $signed(_zz_7730));
  assign _zz_917 = _zz_7731[15 : 0];
  assign _zz_2252 = ($signed(_zz_7732) + $signed(_zz_7733));
  assign _zz_918 = _zz_7734[15 : 0];
  assign _zz_919 = 1'b1;
  assign _zz_920 = 1'b1;
  assign _zz_2253 = ($signed(_zz_7751) - $signed(_zz_7752));
  assign _zz_921 = _zz_7753[15 : 0];
  assign _zz_2254 = ($signed(_zz_7754) + $signed(_zz_7755));
  assign _zz_922 = _zz_7756[15 : 0];
  assign _zz_923 = 1'b1;
  assign _zz_924 = 1'b1;
  assign _zz_2255 = ($signed(_zz_7773) - $signed(_zz_7774));
  assign _zz_925 = _zz_7775[15 : 0];
  assign _zz_2256 = ($signed(_zz_7776) + $signed(_zz_7777));
  assign _zz_926 = _zz_7778[15 : 0];
  assign _zz_927 = 1'b1;
  assign _zz_928 = 1'b1;
  assign _zz_2257 = ($signed(_zz_7795) - $signed(_zz_7796));
  assign _zz_929 = _zz_7797[15 : 0];
  assign _zz_2258 = ($signed(_zz_7798) + $signed(_zz_7799));
  assign _zz_930 = _zz_7800[15 : 0];
  assign _zz_931 = 1'b1;
  assign _zz_932 = 1'b1;
  assign _zz_2259 = ($signed(_zz_7817) - $signed(_zz_7818));
  assign _zz_933 = _zz_7819[15 : 0];
  assign _zz_2260 = ($signed(_zz_7820) + $signed(_zz_7821));
  assign _zz_934 = _zz_7822[15 : 0];
  assign _zz_935 = 1'b1;
  assign _zz_936 = 1'b1;
  assign _zz_2261 = ($signed(_zz_7839) - $signed(_zz_7840));
  assign _zz_937 = _zz_7841[15 : 0];
  assign _zz_2262 = ($signed(_zz_7842) + $signed(_zz_7843));
  assign _zz_938 = _zz_7844[15 : 0];
  assign _zz_939 = 1'b1;
  assign _zz_940 = 1'b1;
  assign _zz_2263 = ($signed(_zz_7861) - $signed(_zz_7862));
  assign _zz_941 = _zz_7863[15 : 0];
  assign _zz_2264 = ($signed(_zz_7864) + $signed(_zz_7865));
  assign _zz_942 = _zz_7866[15 : 0];
  assign _zz_943 = 1'b1;
  assign _zz_944 = 1'b1;
  assign _zz_2265 = ($signed(_zz_7883) - $signed(_zz_7884));
  assign _zz_945 = _zz_7885[15 : 0];
  assign _zz_2266 = ($signed(_zz_7886) + $signed(_zz_7887));
  assign _zz_946 = _zz_7888[15 : 0];
  assign _zz_947 = 1'b1;
  assign _zz_948 = 1'b1;
  assign _zz_2267 = ($signed(_zz_7905) - $signed(_zz_7906));
  assign _zz_949 = _zz_7907[15 : 0];
  assign _zz_2268 = ($signed(_zz_7908) + $signed(_zz_7909));
  assign _zz_950 = _zz_7910[15 : 0];
  assign _zz_951 = 1'b1;
  assign _zz_952 = 1'b1;
  assign _zz_2269 = ($signed(_zz_7927) - $signed(_zz_7928));
  assign _zz_953 = _zz_7929[15 : 0];
  assign _zz_2270 = ($signed(_zz_7930) + $signed(_zz_7931));
  assign _zz_954 = _zz_7932[15 : 0];
  assign _zz_955 = 1'b1;
  assign _zz_956 = 1'b1;
  assign _zz_2271 = ($signed(_zz_7949) - $signed(_zz_7950));
  assign _zz_957 = _zz_7951[15 : 0];
  assign _zz_2272 = ($signed(_zz_7952) + $signed(_zz_7953));
  assign _zz_958 = _zz_7954[15 : 0];
  assign _zz_959 = 1'b1;
  assign _zz_960 = 1'b1;
  assign _zz_2273 = ($signed(_zz_7971) - $signed(_zz_7972));
  assign _zz_961 = _zz_7973[15 : 0];
  assign _zz_2274 = ($signed(_zz_7974) + $signed(_zz_7975));
  assign _zz_962 = _zz_7976[15 : 0];
  assign _zz_963 = 1'b1;
  assign _zz_964 = 1'b1;
  assign _zz_2275 = ($signed(_zz_7993) - $signed(_zz_7994));
  assign _zz_965 = _zz_7995[15 : 0];
  assign _zz_2276 = ($signed(_zz_7996) + $signed(_zz_7997));
  assign _zz_966 = _zz_7998[15 : 0];
  assign _zz_967 = 1'b1;
  assign _zz_968 = 1'b1;
  assign _zz_2277 = ($signed(_zz_8015) - $signed(_zz_8016));
  assign _zz_969 = _zz_8017[15 : 0];
  assign _zz_2278 = ($signed(_zz_8018) + $signed(_zz_8019));
  assign _zz_970 = _zz_8020[15 : 0];
  assign _zz_971 = 1'b1;
  assign _zz_972 = 1'b1;
  assign _zz_2279 = ($signed(_zz_8037) - $signed(_zz_8038));
  assign _zz_973 = _zz_8039[15 : 0];
  assign _zz_2280 = ($signed(_zz_8040) + $signed(_zz_8041));
  assign _zz_974 = _zz_8042[15 : 0];
  assign _zz_975 = 1'b1;
  assign _zz_976 = 1'b1;
  assign _zz_2281 = ($signed(_zz_8059) - $signed(_zz_8060));
  assign _zz_977 = _zz_8061[15 : 0];
  assign _zz_2282 = ($signed(_zz_8062) + $signed(_zz_8063));
  assign _zz_978 = _zz_8064[15 : 0];
  assign _zz_979 = 1'b1;
  assign _zz_980 = 1'b1;
  assign _zz_2283 = ($signed(_zz_8081) - $signed(_zz_8082));
  assign _zz_981 = _zz_8083[15 : 0];
  assign _zz_2284 = ($signed(_zz_8084) + $signed(_zz_8085));
  assign _zz_982 = _zz_8086[15 : 0];
  assign _zz_983 = 1'b1;
  assign _zz_984 = 1'b1;
  assign _zz_2285 = ($signed(_zz_8103) - $signed(_zz_8104));
  assign _zz_985 = _zz_8105[15 : 0];
  assign _zz_2286 = ($signed(_zz_8106) + $signed(_zz_8107));
  assign _zz_986 = _zz_8108[15 : 0];
  assign _zz_987 = 1'b1;
  assign _zz_988 = 1'b1;
  assign _zz_2287 = ($signed(_zz_8125) - $signed(_zz_8126));
  assign _zz_989 = _zz_8127[15 : 0];
  assign _zz_2288 = ($signed(_zz_8128) + $signed(_zz_8129));
  assign _zz_990 = _zz_8130[15 : 0];
  assign _zz_991 = 1'b1;
  assign _zz_992 = 1'b1;
  assign _zz_2289 = ($signed(_zz_8147) - $signed(_zz_8148));
  assign _zz_993 = _zz_8149[15 : 0];
  assign _zz_2290 = ($signed(_zz_8150) + $signed(_zz_8151));
  assign _zz_994 = _zz_8152[15 : 0];
  assign _zz_995 = 1'b1;
  assign _zz_996 = 1'b1;
  assign _zz_2291 = ($signed(_zz_8169) - $signed(_zz_8170));
  assign _zz_997 = _zz_8171[15 : 0];
  assign _zz_2292 = ($signed(_zz_8172) + $signed(_zz_8173));
  assign _zz_998 = _zz_8174[15 : 0];
  assign _zz_999 = 1'b1;
  assign _zz_1000 = 1'b1;
  assign _zz_2293 = ($signed(_zz_8191) - $signed(_zz_8192));
  assign _zz_1001 = _zz_8193[15 : 0];
  assign _zz_2294 = ($signed(_zz_8194) + $signed(_zz_8195));
  assign _zz_1002 = _zz_8196[15 : 0];
  assign _zz_1003 = 1'b1;
  assign _zz_1004 = 1'b1;
  assign _zz_2295 = ($signed(_zz_8213) - $signed(_zz_8214));
  assign _zz_1005 = _zz_8215[15 : 0];
  assign _zz_2296 = ($signed(_zz_8216) + $signed(_zz_8217));
  assign _zz_1006 = _zz_8218[15 : 0];
  assign _zz_1007 = 1'b1;
  assign _zz_1008 = 1'b1;
  assign _zz_2297 = ($signed(_zz_8235) - $signed(_zz_8236));
  assign _zz_1009 = _zz_8237[15 : 0];
  assign _zz_2298 = ($signed(_zz_8238) + $signed(_zz_8239));
  assign _zz_1010 = _zz_8240[15 : 0];
  assign _zz_1011 = 1'b1;
  assign _zz_1012 = 1'b1;
  assign _zz_2299 = ($signed(_zz_8257) - $signed(_zz_8258));
  assign _zz_1013 = _zz_8259[15 : 0];
  assign _zz_2300 = ($signed(_zz_8260) + $signed(_zz_8261));
  assign _zz_1014 = _zz_8262[15 : 0];
  assign _zz_1015 = 1'b1;
  assign _zz_1016 = 1'b1;
  assign _zz_2301 = ($signed(_zz_8279) - $signed(_zz_8280));
  assign _zz_1017 = _zz_8281[15 : 0];
  assign _zz_2302 = ($signed(_zz_8282) + $signed(_zz_8283));
  assign _zz_1018 = _zz_8284[15 : 0];
  assign _zz_1019 = 1'b1;
  assign _zz_1020 = 1'b1;
  assign _zz_2303 = ($signed(_zz_8301) - $signed(_zz_8302));
  assign _zz_1021 = _zz_8303[15 : 0];
  assign _zz_2304 = ($signed(_zz_8304) + $signed(_zz_8305));
  assign _zz_1022 = _zz_8306[15 : 0];
  assign _zz_1023 = 1'b1;
  assign _zz_1024 = 1'b1;
  assign _zz_2305 = ($signed(_zz_8323) - $signed(_zz_8324));
  assign _zz_1025 = _zz_8325[15 : 0];
  assign _zz_2306 = ($signed(_zz_8326) + $signed(_zz_8327));
  assign _zz_1026 = _zz_8328[15 : 0];
  assign _zz_1027 = 1'b1;
  assign _zz_1028 = 1'b1;
  assign _zz_2307 = ($signed(_zz_8345) - $signed(_zz_8346));
  assign _zz_1029 = _zz_8347[15 : 0];
  assign _zz_2308 = ($signed(_zz_8348) + $signed(_zz_8349));
  assign _zz_1030 = _zz_8350[15 : 0];
  assign _zz_1031 = 1'b1;
  assign _zz_1032 = 1'b1;
  assign _zz_2309 = ($signed(_zz_8367) - $signed(_zz_8368));
  assign _zz_1033 = _zz_8369[15 : 0];
  assign _zz_2310 = ($signed(_zz_8370) + $signed(_zz_8371));
  assign _zz_1034 = _zz_8372[15 : 0];
  assign _zz_1035 = 1'b1;
  assign _zz_1036 = 1'b1;
  assign _zz_2311 = ($signed(_zz_8389) - $signed(_zz_8390));
  assign _zz_1037 = _zz_8391[15 : 0];
  assign _zz_2312 = ($signed(_zz_8392) + $signed(_zz_8393));
  assign _zz_1038 = _zz_8394[15 : 0];
  assign _zz_1039 = 1'b1;
  assign _zz_1040 = 1'b1;
  assign _zz_2313 = ($signed(_zz_8411) - $signed(_zz_8412));
  assign _zz_1041 = _zz_8413[15 : 0];
  assign _zz_2314 = ($signed(_zz_8414) + $signed(_zz_8415));
  assign _zz_1042 = _zz_8416[15 : 0];
  assign _zz_1043 = 1'b1;
  assign _zz_1044 = 1'b1;
  assign _zz_2315 = ($signed(_zz_8433) - $signed(_zz_8434));
  assign _zz_1045 = _zz_8435[15 : 0];
  assign _zz_2316 = ($signed(_zz_8436) + $signed(_zz_8437));
  assign _zz_1046 = _zz_8438[15 : 0];
  assign _zz_1047 = 1'b1;
  assign _zz_1048 = 1'b1;
  assign _zz_2317 = ($signed(_zz_8455) - $signed(_zz_8456));
  assign _zz_1049 = _zz_8457[15 : 0];
  assign _zz_2318 = ($signed(_zz_8458) + $signed(_zz_8459));
  assign _zz_1050 = _zz_8460[15 : 0];
  assign _zz_1051 = 1'b1;
  assign _zz_1052 = 1'b1;
  assign _zz_2319 = ($signed(_zz_8477) - $signed(_zz_8478));
  assign _zz_1053 = _zz_8479[15 : 0];
  assign _zz_2320 = ($signed(_zz_8480) + $signed(_zz_8481));
  assign _zz_1054 = _zz_8482[15 : 0];
  assign _zz_1055 = 1'b1;
  assign _zz_1056 = 1'b1;
  assign _zz_2321 = ($signed(_zz_8499) - $signed(_zz_8500));
  assign _zz_1057 = _zz_8501[15 : 0];
  assign _zz_2322 = ($signed(_zz_8502) + $signed(_zz_8503));
  assign _zz_1058 = _zz_8504[15 : 0];
  assign _zz_1059 = 1'b1;
  assign _zz_1060 = 1'b1;
  assign _zz_2323 = ($signed(_zz_8521) - $signed(_zz_8522));
  assign _zz_1061 = _zz_8523[15 : 0];
  assign _zz_2324 = ($signed(_zz_8524) + $signed(_zz_8525));
  assign _zz_1062 = _zz_8526[15 : 0];
  assign _zz_1063 = 1'b1;
  assign _zz_1064 = 1'b1;
  assign _zz_2325 = ($signed(_zz_8543) - $signed(_zz_8544));
  assign _zz_1065 = _zz_8545[15 : 0];
  assign _zz_2326 = ($signed(_zz_8546) + $signed(_zz_8547));
  assign _zz_1066 = _zz_8548[15 : 0];
  assign _zz_1067 = 1'b1;
  assign _zz_1068 = 1'b1;
  assign _zz_2327 = ($signed(_zz_8565) - $signed(_zz_8566));
  assign _zz_1069 = _zz_8567[15 : 0];
  assign _zz_2328 = ($signed(_zz_8568) + $signed(_zz_8569));
  assign _zz_1070 = _zz_8570[15 : 0];
  assign _zz_1071 = 1'b1;
  assign _zz_1072 = 1'b1;
  assign _zz_2329 = ($signed(_zz_8587) - $signed(_zz_8588));
  assign _zz_1073 = _zz_8589[15 : 0];
  assign _zz_2330 = ($signed(_zz_8590) + $signed(_zz_8591));
  assign _zz_1074 = _zz_8592[15 : 0];
  assign _zz_1075 = 1'b1;
  assign _zz_1076 = 1'b1;
  assign _zz_2331 = ($signed(_zz_8609) - $signed(_zz_8610));
  assign _zz_1077 = _zz_8611[15 : 0];
  assign _zz_2332 = ($signed(_zz_8612) + $signed(_zz_8613));
  assign _zz_1078 = _zz_8614[15 : 0];
  assign _zz_1079 = 1'b1;
  assign _zz_1080 = 1'b1;
  assign _zz_2333 = ($signed(_zz_8631) - $signed(_zz_8632));
  assign _zz_1081 = _zz_8633[15 : 0];
  assign _zz_2334 = ($signed(_zz_8634) + $signed(_zz_8635));
  assign _zz_1082 = _zz_8636[15 : 0];
  assign _zz_1083 = 1'b1;
  assign _zz_1084 = 1'b1;
  assign _zz_2335 = ($signed(_zz_8653) - $signed(_zz_8654));
  assign _zz_1085 = _zz_8655[15 : 0];
  assign _zz_2336 = ($signed(_zz_8656) + $signed(_zz_8657));
  assign _zz_1086 = _zz_8658[15 : 0];
  assign _zz_1087 = 1'b1;
  assign _zz_1088 = 1'b1;
  assign _zz_2337 = ($signed(_zz_8675) - $signed(_zz_8676));
  assign _zz_1089 = _zz_8677[15 : 0];
  assign _zz_2338 = ($signed(_zz_8678) + $signed(_zz_8679));
  assign _zz_1090 = _zz_8680[15 : 0];
  assign _zz_1091 = 1'b1;
  assign _zz_1092 = 1'b1;
  assign _zz_2339 = ($signed(_zz_8697) - $signed(_zz_8698));
  assign _zz_1093 = _zz_8699[15 : 0];
  assign _zz_2340 = ($signed(_zz_8700) + $signed(_zz_8701));
  assign _zz_1094 = _zz_8702[15 : 0];
  assign _zz_1095 = 1'b1;
  assign _zz_1096 = 1'b1;
  assign _zz_2341 = ($signed(_zz_8719) - $signed(_zz_8720));
  assign _zz_1097 = _zz_8721[15 : 0];
  assign _zz_2342 = ($signed(_zz_8722) + $signed(_zz_8723));
  assign _zz_1098 = _zz_8724[15 : 0];
  assign _zz_1099 = 1'b1;
  assign _zz_1100 = 1'b1;
  assign _zz_2343 = ($signed(_zz_8741) - $signed(_zz_8742));
  assign _zz_1101 = _zz_8743[15 : 0];
  assign _zz_2344 = ($signed(_zz_8744) + $signed(_zz_8745));
  assign _zz_1102 = _zz_8746[15 : 0];
  assign _zz_1103 = 1'b1;
  assign _zz_1104 = 1'b1;
  assign _zz_2345 = ($signed(_zz_8763) - $signed(_zz_8764));
  assign _zz_1105 = _zz_8765[15 : 0];
  assign _zz_2346 = ($signed(_zz_8766) + $signed(_zz_8767));
  assign _zz_1106 = _zz_8768[15 : 0];
  assign _zz_1107 = 1'b1;
  assign _zz_1108 = 1'b1;
  assign _zz_2347 = ($signed(_zz_8785) - $signed(_zz_8786));
  assign _zz_1109 = _zz_8787[15 : 0];
  assign _zz_2348 = ($signed(_zz_8788) + $signed(_zz_8789));
  assign _zz_1110 = _zz_8790[15 : 0];
  assign _zz_1111 = 1'b1;
  assign _zz_1112 = 1'b1;
  assign _zz_2349 = ($signed(_zz_8807) - $signed(_zz_8808));
  assign _zz_1113 = _zz_8809[15 : 0];
  assign _zz_2350 = ($signed(_zz_8810) + $signed(_zz_8811));
  assign _zz_1114 = _zz_8812[15 : 0];
  assign _zz_1115 = 1'b1;
  assign _zz_1116 = 1'b1;
  assign _zz_2351 = ($signed(_zz_8829) - $signed(_zz_8830));
  assign _zz_1117 = _zz_8831[15 : 0];
  assign _zz_2352 = ($signed(_zz_8832) + $signed(_zz_8833));
  assign _zz_1118 = _zz_8834[15 : 0];
  assign _zz_1119 = 1'b1;
  assign _zz_1120 = 1'b1;
  assign _zz_2353 = ($signed(_zz_8851) - $signed(_zz_8852));
  assign _zz_1121 = _zz_8853[15 : 0];
  assign _zz_2354 = ($signed(_zz_8854) + $signed(_zz_8855));
  assign _zz_1122 = _zz_8856[15 : 0];
  assign _zz_1123 = 1'b1;
  assign _zz_1124 = 1'b1;
  assign _zz_2355 = ($signed(_zz_8873) - $signed(_zz_8874));
  assign _zz_1125 = _zz_8875[15 : 0];
  assign _zz_2356 = ($signed(_zz_8876) + $signed(_zz_8877));
  assign _zz_1126 = _zz_8878[15 : 0];
  assign _zz_1127 = 1'b1;
  assign _zz_1128 = 1'b1;
  assign _zz_2357 = ($signed(_zz_8895) - $signed(_zz_8896));
  assign _zz_1129 = _zz_8897[15 : 0];
  assign _zz_2358 = ($signed(_zz_8898) + $signed(_zz_8899));
  assign _zz_1130 = _zz_8900[15 : 0];
  assign _zz_1131 = 1'b1;
  assign _zz_1132 = 1'b1;
  assign _zz_2359 = ($signed(_zz_8917) - $signed(_zz_8918));
  assign _zz_1133 = _zz_8919[15 : 0];
  assign _zz_2360 = ($signed(_zz_8920) + $signed(_zz_8921));
  assign _zz_1134 = _zz_8922[15 : 0];
  assign _zz_1135 = 1'b1;
  assign _zz_1136 = 1'b1;
  assign _zz_2361 = ($signed(_zz_8939) - $signed(_zz_8940));
  assign _zz_1137 = _zz_8941[15 : 0];
  assign _zz_2362 = ($signed(_zz_8942) + $signed(_zz_8943));
  assign _zz_1138 = _zz_8944[15 : 0];
  assign _zz_1139 = 1'b1;
  assign _zz_1140 = 1'b1;
  assign _zz_2363 = ($signed(_zz_8961) - $signed(_zz_8962));
  assign _zz_1141 = _zz_8963[15 : 0];
  assign _zz_2364 = ($signed(_zz_8964) + $signed(_zz_8965));
  assign _zz_1142 = _zz_8966[15 : 0];
  assign _zz_1143 = 1'b1;
  assign _zz_1144 = 1'b1;
  assign _zz_2365 = ($signed(_zz_8983) - $signed(_zz_8984));
  assign _zz_1145 = _zz_8985[15 : 0];
  assign _zz_2366 = ($signed(_zz_8986) + $signed(_zz_8987));
  assign _zz_1146 = _zz_8988[15 : 0];
  assign _zz_1147 = 1'b1;
  assign _zz_1148 = 1'b1;
  assign _zz_2367 = ($signed(_zz_9005) - $signed(_zz_9006));
  assign _zz_1149 = _zz_9007[15 : 0];
  assign _zz_2368 = ($signed(_zz_9008) + $signed(_zz_9009));
  assign _zz_1150 = _zz_9010[15 : 0];
  assign _zz_1151 = 1'b1;
  assign _zz_1152 = 1'b1;
  assign _zz_2369 = ($signed(_zz_9027) - $signed(_zz_9028));
  assign _zz_1153 = _zz_9029[15 : 0];
  assign _zz_2370 = ($signed(_zz_9030) + $signed(_zz_9031));
  assign _zz_1154 = _zz_9032[15 : 0];
  assign _zz_1155 = 1'b1;
  assign _zz_1156 = 1'b1;
  assign _zz_2371 = ($signed(_zz_9049) - $signed(_zz_9050));
  assign _zz_1157 = _zz_9051[15 : 0];
  assign _zz_2372 = ($signed(_zz_9052) + $signed(_zz_9053));
  assign _zz_1158 = _zz_9054[15 : 0];
  assign _zz_1159 = 1'b1;
  assign _zz_1160 = 1'b1;
  assign _zz_2373 = ($signed(_zz_9071) - $signed(_zz_9072));
  assign _zz_1161 = _zz_9073[15 : 0];
  assign _zz_2374 = ($signed(_zz_9074) + $signed(_zz_9075));
  assign _zz_1162 = _zz_9076[15 : 0];
  assign _zz_1163 = 1'b1;
  assign _zz_1164 = 1'b1;
  assign _zz_2375 = ($signed(_zz_9093) - $signed(_zz_9094));
  assign _zz_1165 = _zz_9095[15 : 0];
  assign _zz_2376 = ($signed(_zz_9096) + $signed(_zz_9097));
  assign _zz_1166 = _zz_9098[15 : 0];
  assign _zz_1167 = 1'b1;
  assign _zz_1168 = 1'b1;
  assign _zz_2377 = ($signed(_zz_9115) - $signed(_zz_9116));
  assign _zz_1169 = _zz_9117[15 : 0];
  assign _zz_2378 = ($signed(_zz_9118) + $signed(_zz_9119));
  assign _zz_1170 = _zz_9120[15 : 0];
  assign _zz_1171 = 1'b1;
  assign _zz_1172 = 1'b1;
  assign _zz_2379 = ($signed(_zz_9137) - $signed(_zz_9138));
  assign _zz_1173 = _zz_9139[15 : 0];
  assign _zz_2380 = ($signed(_zz_9140) + $signed(_zz_9141));
  assign _zz_1174 = _zz_9142[15 : 0];
  assign _zz_1175 = 1'b1;
  assign _zz_1176 = 1'b1;
  assign _zz_2381 = ($signed(_zz_9159) - $signed(_zz_9160));
  assign _zz_1177 = _zz_9161[15 : 0];
  assign _zz_2382 = ($signed(_zz_9162) + $signed(_zz_9163));
  assign _zz_1178 = _zz_9164[15 : 0];
  assign _zz_1179 = 1'b1;
  assign _zz_1180 = 1'b1;
  assign _zz_2383 = ($signed(_zz_9181) - $signed(_zz_9182));
  assign _zz_1181 = _zz_9183[15 : 0];
  assign _zz_2384 = ($signed(_zz_9184) + $signed(_zz_9185));
  assign _zz_1182 = _zz_9186[15 : 0];
  assign _zz_1183 = 1'b1;
  assign _zz_1184 = 1'b1;
  assign _zz_2385 = ($signed(_zz_9203) - $signed(_zz_9204));
  assign _zz_1185 = _zz_9205[15 : 0];
  assign _zz_2386 = ($signed(_zz_9206) + $signed(_zz_9207));
  assign _zz_1186 = _zz_9208[15 : 0];
  assign _zz_1187 = 1'b1;
  assign _zz_1188 = 1'b1;
  assign _zz_2387 = ($signed(_zz_9225) - $signed(_zz_9226));
  assign _zz_1189 = _zz_9227[15 : 0];
  assign _zz_2388 = ($signed(_zz_9228) + $signed(_zz_9229));
  assign _zz_1190 = _zz_9230[15 : 0];
  assign _zz_1191 = 1'b1;
  assign _zz_1192 = 1'b1;
  assign _zz_2389 = ($signed(_zz_9247) - $signed(_zz_9248));
  assign _zz_1193 = _zz_9249[15 : 0];
  assign _zz_2390 = ($signed(_zz_9250) + $signed(_zz_9251));
  assign _zz_1194 = _zz_9252[15 : 0];
  assign _zz_1195 = 1'b1;
  assign _zz_1196 = 1'b1;
  assign _zz_2391 = ($signed(_zz_9269) - $signed(_zz_9270));
  assign _zz_1197 = _zz_9271[15 : 0];
  assign _zz_2392 = ($signed(_zz_9272) + $signed(_zz_9273));
  assign _zz_1198 = _zz_9274[15 : 0];
  assign _zz_1199 = 1'b1;
  assign _zz_1200 = 1'b1;
  assign _zz_2393 = ($signed(_zz_9291) - $signed(_zz_9292));
  assign _zz_1201 = _zz_9293[15 : 0];
  assign _zz_2394 = ($signed(_zz_9294) + $signed(_zz_9295));
  assign _zz_1202 = _zz_9296[15 : 0];
  assign _zz_1203 = 1'b1;
  assign _zz_1204 = 1'b1;
  assign _zz_2395 = ($signed(_zz_9313) - $signed(_zz_9314));
  assign _zz_1205 = _zz_9315[15 : 0];
  assign _zz_2396 = ($signed(_zz_9316) + $signed(_zz_9317));
  assign _zz_1206 = _zz_9318[15 : 0];
  assign _zz_1207 = 1'b1;
  assign _zz_1208 = 1'b1;
  assign _zz_2397 = ($signed(_zz_9335) - $signed(_zz_9336));
  assign _zz_1209 = _zz_9337[15 : 0];
  assign _zz_2398 = ($signed(_zz_9338) + $signed(_zz_9339));
  assign _zz_1210 = _zz_9340[15 : 0];
  assign _zz_1211 = 1'b1;
  assign _zz_1212 = 1'b1;
  assign _zz_2399 = ($signed(_zz_9357) - $signed(_zz_9358));
  assign _zz_1213 = _zz_9359[15 : 0];
  assign _zz_2400 = ($signed(_zz_9360) + $signed(_zz_9361));
  assign _zz_1214 = _zz_9362[15 : 0];
  assign _zz_1215 = 1'b1;
  assign _zz_1216 = 1'b1;
  assign _zz_2401 = ($signed(_zz_9379) - $signed(_zz_9380));
  assign _zz_1217 = _zz_9381[15 : 0];
  assign _zz_2402 = ($signed(_zz_9382) + $signed(_zz_9383));
  assign _zz_1218 = _zz_9384[15 : 0];
  assign _zz_1219 = 1'b1;
  assign _zz_1220 = 1'b1;
  assign _zz_2403 = ($signed(_zz_9401) - $signed(_zz_9402));
  assign _zz_1221 = _zz_9403[15 : 0];
  assign _zz_2404 = ($signed(_zz_9404) + $signed(_zz_9405));
  assign _zz_1222 = _zz_9406[15 : 0];
  assign _zz_1223 = 1'b1;
  assign _zz_1224 = 1'b1;
  assign _zz_2405 = ($signed(_zz_9423) - $signed(_zz_9424));
  assign _zz_1225 = _zz_9425[15 : 0];
  assign _zz_2406 = ($signed(_zz_9426) + $signed(_zz_9427));
  assign _zz_1226 = _zz_9428[15 : 0];
  assign _zz_1227 = 1'b1;
  assign _zz_1228 = 1'b1;
  assign _zz_2407 = ($signed(_zz_9445) - $signed(_zz_9446));
  assign _zz_1229 = _zz_9447[15 : 0];
  assign _zz_2408 = ($signed(_zz_9448) + $signed(_zz_9449));
  assign _zz_1230 = _zz_9450[15 : 0];
  assign _zz_1231 = 1'b1;
  assign _zz_1232 = 1'b1;
  assign _zz_2409 = ($signed(_zz_9467) - $signed(_zz_9468));
  assign _zz_1233 = _zz_9469[15 : 0];
  assign _zz_2410 = ($signed(_zz_9470) + $signed(_zz_9471));
  assign _zz_1234 = _zz_9472[15 : 0];
  assign _zz_1235 = 1'b1;
  assign _zz_1236 = 1'b1;
  assign _zz_2411 = ($signed(_zz_9489) - $signed(_zz_9490));
  assign _zz_1237 = _zz_9491[15 : 0];
  assign _zz_2412 = ($signed(_zz_9492) + $signed(_zz_9493));
  assign _zz_1238 = _zz_9494[15 : 0];
  assign _zz_1239 = 1'b1;
  assign _zz_1240 = 1'b1;
  assign _zz_2413 = ($signed(_zz_9511) - $signed(_zz_9512));
  assign _zz_1241 = _zz_9513[15 : 0];
  assign _zz_2414 = ($signed(_zz_9514) + $signed(_zz_9515));
  assign _zz_1242 = _zz_9516[15 : 0];
  assign _zz_1243 = 1'b1;
  assign _zz_1244 = 1'b1;
  assign _zz_2415 = ($signed(_zz_9533) - $signed(_zz_9534));
  assign _zz_1245 = _zz_9535[15 : 0];
  assign _zz_2416 = ($signed(_zz_9536) + $signed(_zz_9537));
  assign _zz_1246 = _zz_9538[15 : 0];
  assign _zz_1247 = 1'b1;
  assign _zz_1248 = 1'b1;
  assign _zz_2417 = ($signed(_zz_9555) - $signed(_zz_9556));
  assign _zz_1249 = _zz_9557[15 : 0];
  assign _zz_2418 = ($signed(_zz_9558) + $signed(_zz_9559));
  assign _zz_1250 = _zz_9560[15 : 0];
  assign _zz_1251 = 1'b1;
  assign _zz_1252 = 1'b1;
  assign _zz_2419 = ($signed(_zz_9577) - $signed(_zz_9578));
  assign _zz_1253 = _zz_9579[15 : 0];
  assign _zz_2420 = ($signed(_zz_9580) + $signed(_zz_9581));
  assign _zz_1254 = _zz_9582[15 : 0];
  assign _zz_1255 = 1'b1;
  assign _zz_1256 = 1'b1;
  assign _zz_2421 = ($signed(_zz_9599) - $signed(_zz_9600));
  assign _zz_1257 = _zz_9601[15 : 0];
  assign _zz_2422 = ($signed(_zz_9602) + $signed(_zz_9603));
  assign _zz_1258 = _zz_9604[15 : 0];
  assign _zz_1259 = 1'b1;
  assign _zz_1260 = 1'b1;
  assign _zz_2423 = ($signed(_zz_9621) - $signed(_zz_9622));
  assign _zz_1261 = _zz_9623[15 : 0];
  assign _zz_2424 = ($signed(_zz_9624) + $signed(_zz_9625));
  assign _zz_1262 = _zz_9626[15 : 0];
  assign _zz_1263 = 1'b1;
  assign _zz_1264 = 1'b1;
  assign _zz_2425 = ($signed(_zz_9643) - $signed(_zz_9644));
  assign _zz_1265 = _zz_9645[15 : 0];
  assign _zz_2426 = ($signed(_zz_9646) + $signed(_zz_9647));
  assign _zz_1266 = _zz_9648[15 : 0];
  assign _zz_1267 = 1'b1;
  assign _zz_1268 = 1'b1;
  assign _zz_2427 = ($signed(_zz_9665) - $signed(_zz_9666));
  assign _zz_1269 = _zz_9667[15 : 0];
  assign _zz_2428 = ($signed(_zz_9668) + $signed(_zz_9669));
  assign _zz_1270 = _zz_9670[15 : 0];
  assign _zz_1271 = 1'b1;
  assign _zz_1272 = 1'b1;
  assign _zz_2429 = ($signed(_zz_9687) - $signed(_zz_9688));
  assign _zz_1273 = _zz_9689[15 : 0];
  assign _zz_2430 = ($signed(_zz_9690) + $signed(_zz_9691));
  assign _zz_1274 = _zz_9692[15 : 0];
  assign _zz_1275 = 1'b1;
  assign _zz_1276 = 1'b1;
  assign _zz_2431 = ($signed(_zz_9709) - $signed(_zz_9710));
  assign _zz_1277 = _zz_9711[15 : 0];
  assign _zz_2432 = ($signed(_zz_9712) + $signed(_zz_9713));
  assign _zz_1278 = _zz_9714[15 : 0];
  assign _zz_1279 = 1'b1;
  assign _zz_1280 = 1'b1;
  assign _zz_2433 = ($signed(_zz_9731) - $signed(_zz_9732));
  assign _zz_1281 = _zz_9733[15 : 0];
  assign _zz_2434 = ($signed(_zz_9734) + $signed(_zz_9735));
  assign _zz_1282 = _zz_9736[15 : 0];
  assign _zz_1283 = 1'b1;
  assign _zz_1284 = 1'b1;
  assign _zz_2435 = ($signed(_zz_9753) - $signed(_zz_9754));
  assign _zz_1285 = _zz_9755[15 : 0];
  assign _zz_2436 = ($signed(_zz_9756) + $signed(_zz_9757));
  assign _zz_1286 = _zz_9758[15 : 0];
  assign _zz_1287 = 1'b1;
  assign _zz_1288 = 1'b1;
  assign _zz_2437 = ($signed(_zz_9775) - $signed(_zz_9776));
  assign _zz_1289 = _zz_9777[15 : 0];
  assign _zz_2438 = ($signed(_zz_9778) + $signed(_zz_9779));
  assign _zz_1290 = _zz_9780[15 : 0];
  assign _zz_1291 = 1'b1;
  assign _zz_1292 = 1'b1;
  assign _zz_2439 = ($signed(_zz_9797) - $signed(_zz_9798));
  assign _zz_1293 = _zz_9799[15 : 0];
  assign _zz_2440 = ($signed(_zz_9800) + $signed(_zz_9801));
  assign _zz_1294 = _zz_9802[15 : 0];
  assign _zz_1295 = 1'b1;
  assign _zz_1296 = 1'b1;
  assign _zz_2441 = ($signed(_zz_9819) - $signed(_zz_9820));
  assign _zz_1297 = _zz_9821[15 : 0];
  assign _zz_2442 = ($signed(_zz_9822) + $signed(_zz_9823));
  assign _zz_1298 = _zz_9824[15 : 0];
  assign _zz_1299 = 1'b1;
  assign _zz_1300 = 1'b1;
  assign _zz_2443 = ($signed(_zz_9841) - $signed(_zz_9842));
  assign _zz_1301 = _zz_9843[15 : 0];
  assign _zz_2444 = ($signed(_zz_9844) + $signed(_zz_9845));
  assign _zz_1302 = _zz_9846[15 : 0];
  assign _zz_1303 = 1'b1;
  assign _zz_1304 = 1'b1;
  assign _zz_2445 = ($signed(_zz_9863) - $signed(_zz_9864));
  assign _zz_1305 = _zz_9865[15 : 0];
  assign _zz_2446 = ($signed(_zz_9866) + $signed(_zz_9867));
  assign _zz_1306 = _zz_9868[15 : 0];
  assign _zz_1307 = 1'b1;
  assign _zz_1308 = 1'b1;
  assign _zz_2447 = ($signed(_zz_9885) - $signed(_zz_9886));
  assign _zz_1309 = _zz_9887[15 : 0];
  assign _zz_2448 = ($signed(_zz_9888) + $signed(_zz_9889));
  assign _zz_1310 = _zz_9890[15 : 0];
  assign _zz_1311 = 1'b1;
  assign _zz_1312 = 1'b1;
  assign _zz_2449 = ($signed(_zz_9907) - $signed(_zz_9908));
  assign _zz_1313 = _zz_9909[15 : 0];
  assign _zz_2450 = ($signed(_zz_9910) + $signed(_zz_9911));
  assign _zz_1314 = _zz_9912[15 : 0];
  assign _zz_1315 = 1'b1;
  assign _zz_1316 = 1'b1;
  assign _zz_2451 = ($signed(_zz_9929) - $signed(_zz_9930));
  assign _zz_1317 = _zz_9931[15 : 0];
  assign _zz_2452 = ($signed(_zz_9932) + $signed(_zz_9933));
  assign _zz_1318 = _zz_9934[15 : 0];
  assign _zz_1319 = 1'b1;
  assign _zz_1320 = 1'b1;
  assign _zz_2453 = ($signed(_zz_9951) - $signed(_zz_9952));
  assign _zz_1321 = _zz_9953[15 : 0];
  assign _zz_2454 = ($signed(_zz_9954) + $signed(_zz_9955));
  assign _zz_1322 = _zz_9956[15 : 0];
  assign _zz_1323 = 1'b1;
  assign _zz_1324 = 1'b1;
  assign _zz_2455 = ($signed(_zz_9973) - $signed(_zz_9974));
  assign _zz_1325 = _zz_9975[15 : 0];
  assign _zz_2456 = ($signed(_zz_9976) + $signed(_zz_9977));
  assign _zz_1326 = _zz_9978[15 : 0];
  assign _zz_1327 = 1'b1;
  assign _zz_1328 = 1'b1;
  assign _zz_2457 = ($signed(_zz_9995) - $signed(_zz_9996));
  assign _zz_1329 = _zz_9997[15 : 0];
  assign _zz_2458 = ($signed(_zz_9998) + $signed(_zz_9999));
  assign _zz_1330 = _zz_10000[15 : 0];
  assign _zz_1331 = 1'b1;
  assign _zz_1332 = 1'b1;
  assign _zz_2459 = ($signed(_zz_10017) - $signed(_zz_10018));
  assign _zz_1333 = _zz_10019[15 : 0];
  assign _zz_2460 = ($signed(_zz_10020) + $signed(_zz_10021));
  assign _zz_1334 = _zz_10022[15 : 0];
  assign _zz_1335 = 1'b1;
  assign _zz_1336 = 1'b1;
  assign _zz_2461 = ($signed(_zz_10039) - $signed(_zz_10040));
  assign _zz_1337 = _zz_10041[15 : 0];
  assign _zz_2462 = ($signed(_zz_10042) + $signed(_zz_10043));
  assign _zz_1338 = _zz_10044[15 : 0];
  assign _zz_1339 = 1'b1;
  assign _zz_1340 = 1'b1;
  assign _zz_2463 = ($signed(_zz_10061) - $signed(_zz_10062));
  assign _zz_1341 = _zz_10063[15 : 0];
  assign _zz_2464 = ($signed(_zz_10064) + $signed(_zz_10065));
  assign _zz_1342 = _zz_10066[15 : 0];
  assign _zz_1343 = 1'b1;
  assign _zz_1344 = 1'b1;
  assign _zz_2465 = ($signed(_zz_10083) - $signed(_zz_10084));
  assign _zz_1345 = _zz_10085[15 : 0];
  assign _zz_2466 = ($signed(_zz_10086) + $signed(_zz_10087));
  assign _zz_1346 = _zz_10088[15 : 0];
  assign _zz_1347 = 1'b1;
  assign _zz_1348 = 1'b1;
  assign _zz_2467 = ($signed(_zz_10105) - $signed(_zz_10106));
  assign _zz_1349 = _zz_10107[15 : 0];
  assign _zz_2468 = ($signed(_zz_10108) + $signed(_zz_10109));
  assign _zz_1350 = _zz_10110[15 : 0];
  assign _zz_1351 = 1'b1;
  assign _zz_1352 = 1'b1;
  assign _zz_2469 = ($signed(_zz_10127) - $signed(_zz_10128));
  assign _zz_1353 = _zz_10129[15 : 0];
  assign _zz_2470 = ($signed(_zz_10130) + $signed(_zz_10131));
  assign _zz_1354 = _zz_10132[15 : 0];
  assign _zz_1355 = 1'b1;
  assign _zz_1356 = 1'b1;
  assign _zz_2471 = ($signed(_zz_10149) - $signed(_zz_10150));
  assign _zz_1357 = _zz_10151[15 : 0];
  assign _zz_2472 = ($signed(_zz_10152) + $signed(_zz_10153));
  assign _zz_1358 = _zz_10154[15 : 0];
  assign _zz_1359 = 1'b1;
  assign _zz_1360 = 1'b1;
  assign _zz_2473 = ($signed(_zz_10171) - $signed(_zz_10172));
  assign _zz_1361 = _zz_10173[15 : 0];
  assign _zz_2474 = ($signed(_zz_10174) + $signed(_zz_10175));
  assign _zz_1362 = _zz_10176[15 : 0];
  assign _zz_1363 = 1'b1;
  assign _zz_1364 = 1'b1;
  assign _zz_2475 = ($signed(_zz_10193) - $signed(_zz_10194));
  assign _zz_1365 = _zz_10195[15 : 0];
  assign _zz_2476 = ($signed(_zz_10196) + $signed(_zz_10197));
  assign _zz_1366 = _zz_10198[15 : 0];
  assign _zz_1367 = 1'b1;
  assign _zz_1368 = 1'b1;
  assign _zz_2477 = ($signed(_zz_10215) - $signed(_zz_10216));
  assign _zz_1369 = _zz_10217[15 : 0];
  assign _zz_2478 = ($signed(_zz_10218) + $signed(_zz_10219));
  assign _zz_1370 = _zz_10220[15 : 0];
  assign _zz_1371 = 1'b1;
  assign _zz_1372 = 1'b1;
  assign _zz_2479 = ($signed(_zz_10237) - $signed(_zz_10238));
  assign _zz_1373 = _zz_10239[15 : 0];
  assign _zz_2480 = ($signed(_zz_10240) + $signed(_zz_10241));
  assign _zz_1374 = _zz_10242[15 : 0];
  assign _zz_1375 = 1'b1;
  assign _zz_1376 = 1'b1;
  assign _zz_2481 = ($signed(_zz_10259) - $signed(_zz_10260));
  assign _zz_1377 = _zz_10261[15 : 0];
  assign _zz_2482 = ($signed(_zz_10262) + $signed(_zz_10263));
  assign _zz_1378 = _zz_10264[15 : 0];
  assign _zz_1379 = 1'b1;
  assign _zz_1380 = 1'b1;
  assign _zz_2483 = ($signed(_zz_10281) - $signed(_zz_10282));
  assign _zz_1381 = _zz_10283[15 : 0];
  assign _zz_2484 = ($signed(_zz_10284) + $signed(_zz_10285));
  assign _zz_1382 = _zz_10286[15 : 0];
  assign _zz_1383 = 1'b1;
  assign _zz_1384 = 1'b1;
  assign _zz_2485 = ($signed(_zz_10303) - $signed(_zz_10304));
  assign _zz_1385 = _zz_10305[15 : 0];
  assign _zz_2486 = ($signed(_zz_10306) + $signed(_zz_10307));
  assign _zz_1386 = _zz_10308[15 : 0];
  assign _zz_1387 = 1'b1;
  assign _zz_1388 = 1'b1;
  assign _zz_2487 = ($signed(_zz_10325) - $signed(_zz_10326));
  assign _zz_1389 = _zz_10327[15 : 0];
  assign _zz_2488 = ($signed(_zz_10328) + $signed(_zz_10329));
  assign _zz_1390 = _zz_10330[15 : 0];
  assign _zz_1391 = 1'b1;
  assign _zz_1392 = 1'b1;
  assign _zz_2489 = ($signed(_zz_10347) - $signed(_zz_10348));
  assign _zz_1393 = _zz_10349[15 : 0];
  assign _zz_2490 = ($signed(_zz_10350) + $signed(_zz_10351));
  assign _zz_1394 = _zz_10352[15 : 0];
  assign _zz_1395 = 1'b1;
  assign _zz_1396 = 1'b1;
  assign _zz_2491 = ($signed(_zz_10369) - $signed(_zz_10370));
  assign _zz_1397 = _zz_10371[15 : 0];
  assign _zz_2492 = ($signed(_zz_10372) + $signed(_zz_10373));
  assign _zz_1398 = _zz_10374[15 : 0];
  assign _zz_1399 = 1'b1;
  assign _zz_1400 = 1'b1;
  assign _zz_2493 = ($signed(_zz_10391) - $signed(_zz_10392));
  assign _zz_1401 = _zz_10393[15 : 0];
  assign _zz_2494 = ($signed(_zz_10394) + $signed(_zz_10395));
  assign _zz_1402 = _zz_10396[15 : 0];
  assign _zz_1403 = 1'b1;
  assign _zz_1404 = 1'b1;
  assign _zz_2495 = ($signed(_zz_10413) - $signed(_zz_10414));
  assign _zz_1405 = _zz_10415[15 : 0];
  assign _zz_2496 = ($signed(_zz_10416) + $signed(_zz_10417));
  assign _zz_1406 = _zz_10418[15 : 0];
  assign _zz_1407 = 1'b1;
  assign _zz_1408 = 1'b1;
  assign _zz_2497 = ($signed(_zz_10435) - $signed(_zz_10436));
  assign _zz_1409 = _zz_10437[15 : 0];
  assign _zz_2498 = ($signed(_zz_10438) + $signed(_zz_10439));
  assign _zz_1410 = _zz_10440[15 : 0];
  assign _zz_1411 = 1'b1;
  assign _zz_1412 = 1'b1;
  assign _zz_2499 = ($signed(_zz_10457) - $signed(_zz_10458));
  assign _zz_1413 = _zz_10459[15 : 0];
  assign _zz_2500 = ($signed(_zz_10460) + $signed(_zz_10461));
  assign _zz_1414 = _zz_10462[15 : 0];
  assign _zz_1415 = 1'b1;
  assign _zz_1416 = 1'b1;
  assign _zz_2501 = ($signed(_zz_10479) - $signed(_zz_10480));
  assign _zz_1417 = _zz_10481[15 : 0];
  assign _zz_2502 = ($signed(_zz_10482) + $signed(_zz_10483));
  assign _zz_1418 = _zz_10484[15 : 0];
  assign _zz_1419 = 1'b1;
  assign _zz_1420 = 1'b1;
  assign _zz_2503 = ($signed(_zz_10501) - $signed(_zz_10502));
  assign _zz_1421 = _zz_10503[15 : 0];
  assign _zz_2504 = ($signed(_zz_10504) + $signed(_zz_10505));
  assign _zz_1422 = _zz_10506[15 : 0];
  assign _zz_1423 = 1'b1;
  assign _zz_1424 = 1'b1;
  assign _zz_2505 = ($signed(_zz_10523) - $signed(_zz_10524));
  assign _zz_1425 = _zz_10525[15 : 0];
  assign _zz_2506 = ($signed(_zz_10526) + $signed(_zz_10527));
  assign _zz_1426 = _zz_10528[15 : 0];
  assign _zz_1427 = 1'b1;
  assign _zz_1428 = 1'b1;
  assign _zz_2507 = ($signed(_zz_10545) - $signed(_zz_10546));
  assign _zz_1429 = _zz_10547[15 : 0];
  assign _zz_2508 = ($signed(_zz_10548) + $signed(_zz_10549));
  assign _zz_1430 = _zz_10550[15 : 0];
  assign _zz_1431 = 1'b1;
  assign _zz_1432 = 1'b1;
  assign _zz_2509 = ($signed(_zz_10567) - $signed(_zz_10568));
  assign _zz_1433 = _zz_10569[15 : 0];
  assign _zz_2510 = ($signed(_zz_10570) + $signed(_zz_10571));
  assign _zz_1434 = _zz_10572[15 : 0];
  assign _zz_1435 = 1'b1;
  assign _zz_1436 = 1'b1;
  assign _zz_2511 = ($signed(_zz_10589) - $signed(_zz_10590));
  assign _zz_1437 = _zz_10591[15 : 0];
  assign _zz_2512 = ($signed(_zz_10592) + $signed(_zz_10593));
  assign _zz_1438 = _zz_10594[15 : 0];
  assign _zz_1439 = 1'b1;
  assign _zz_1440 = 1'b1;
  assign _zz_2513 = ($signed(_zz_10611) - $signed(_zz_10612));
  assign _zz_1441 = _zz_10613[15 : 0];
  assign _zz_2514 = ($signed(_zz_10614) + $signed(_zz_10615));
  assign _zz_1442 = _zz_10616[15 : 0];
  assign _zz_1443 = 1'b1;
  assign _zz_1444 = 1'b1;
  assign _zz_2515 = ($signed(_zz_10633) - $signed(_zz_10634));
  assign _zz_1445 = _zz_10635[15 : 0];
  assign _zz_2516 = ($signed(_zz_10636) + $signed(_zz_10637));
  assign _zz_1446 = _zz_10638[15 : 0];
  assign _zz_1447 = 1'b1;
  assign _zz_1448 = 1'b1;
  assign _zz_2517 = ($signed(_zz_10655) - $signed(_zz_10656));
  assign _zz_1449 = _zz_10657[15 : 0];
  assign _zz_2518 = ($signed(_zz_10658) + $signed(_zz_10659));
  assign _zz_1450 = _zz_10660[15 : 0];
  assign _zz_1451 = 1'b1;
  assign _zz_1452 = 1'b1;
  assign _zz_2519 = ($signed(_zz_10677) - $signed(_zz_10678));
  assign _zz_1453 = _zz_10679[15 : 0];
  assign _zz_2520 = ($signed(_zz_10680) + $signed(_zz_10681));
  assign _zz_1454 = _zz_10682[15 : 0];
  assign _zz_1455 = 1'b1;
  assign _zz_1456 = 1'b1;
  assign _zz_2521 = ($signed(_zz_10699) - $signed(_zz_10700));
  assign _zz_1457 = _zz_10701[15 : 0];
  assign _zz_2522 = ($signed(_zz_10702) + $signed(_zz_10703));
  assign _zz_1458 = _zz_10704[15 : 0];
  assign _zz_1459 = 1'b1;
  assign _zz_1460 = 1'b1;
  assign _zz_2523 = ($signed(_zz_10721) - $signed(_zz_10722));
  assign _zz_1461 = _zz_10723[15 : 0];
  assign _zz_2524 = ($signed(_zz_10724) + $signed(_zz_10725));
  assign _zz_1462 = _zz_10726[15 : 0];
  assign _zz_1463 = 1'b1;
  assign _zz_1464 = 1'b1;
  assign _zz_2525 = ($signed(_zz_10743) - $signed(_zz_10744));
  assign _zz_1465 = _zz_10745[15 : 0];
  assign _zz_2526 = ($signed(_zz_10746) + $signed(_zz_10747));
  assign _zz_1466 = _zz_10748[15 : 0];
  assign _zz_1467 = 1'b1;
  assign _zz_1468 = 1'b1;
  assign _zz_2527 = ($signed(_zz_10765) - $signed(_zz_10766));
  assign _zz_1469 = _zz_10767[15 : 0];
  assign _zz_2528 = ($signed(_zz_10768) + $signed(_zz_10769));
  assign _zz_1470 = _zz_10770[15 : 0];
  assign _zz_1471 = 1'b1;
  assign _zz_1472 = 1'b1;
  assign _zz_2529 = ($signed(_zz_10787) - $signed(_zz_10788));
  assign _zz_1473 = _zz_10789[15 : 0];
  assign _zz_2530 = ($signed(_zz_10790) + $signed(_zz_10791));
  assign _zz_1474 = _zz_10792[15 : 0];
  assign _zz_1475 = 1'b1;
  assign _zz_1476 = 1'b1;
  assign _zz_2531 = ($signed(_zz_10809) - $signed(_zz_10810));
  assign _zz_1477 = _zz_10811[15 : 0];
  assign _zz_2532 = ($signed(_zz_10812) + $signed(_zz_10813));
  assign _zz_1478 = _zz_10814[15 : 0];
  assign _zz_1479 = 1'b1;
  assign _zz_1480 = 1'b1;
  assign _zz_2533 = ($signed(_zz_10831) - $signed(_zz_10832));
  assign _zz_1481 = _zz_10833[15 : 0];
  assign _zz_2534 = ($signed(_zz_10834) + $signed(_zz_10835));
  assign _zz_1482 = _zz_10836[15 : 0];
  assign _zz_1483 = 1'b1;
  assign _zz_1484 = 1'b1;
  assign _zz_2535 = ($signed(_zz_10853) - $signed(_zz_10854));
  assign _zz_1485 = _zz_10855[15 : 0];
  assign _zz_2536 = ($signed(_zz_10856) + $signed(_zz_10857));
  assign _zz_1486 = _zz_10858[15 : 0];
  assign _zz_1487 = 1'b1;
  assign _zz_1488 = 1'b1;
  assign _zz_2537 = ($signed(_zz_10875) - $signed(_zz_10876));
  assign _zz_1489 = _zz_10877[15 : 0];
  assign _zz_2538 = ($signed(_zz_10878) + $signed(_zz_10879));
  assign _zz_1490 = _zz_10880[15 : 0];
  assign _zz_1491 = 1'b1;
  assign _zz_1492 = 1'b1;
  assign _zz_2539 = ($signed(_zz_10897) - $signed(_zz_10898));
  assign _zz_1493 = _zz_10899[15 : 0];
  assign _zz_2540 = ($signed(_zz_10900) + $signed(_zz_10901));
  assign _zz_1494 = _zz_10902[15 : 0];
  assign _zz_1495 = 1'b1;
  assign _zz_1496 = 1'b1;
  assign _zz_2541 = ($signed(_zz_10919) - $signed(_zz_10920));
  assign _zz_1497 = _zz_10921[15 : 0];
  assign _zz_2542 = ($signed(_zz_10922) + $signed(_zz_10923));
  assign _zz_1498 = _zz_10924[15 : 0];
  assign _zz_1499 = 1'b1;
  assign _zz_1500 = 1'b1;
  assign _zz_2543 = ($signed(_zz_10941) - $signed(_zz_10942));
  assign _zz_1501 = _zz_10943[15 : 0];
  assign _zz_2544 = ($signed(_zz_10944) + $signed(_zz_10945));
  assign _zz_1502 = _zz_10946[15 : 0];
  assign _zz_1503 = 1'b1;
  assign _zz_1504 = 1'b1;
  assign _zz_2545 = ($signed(_zz_10963) - $signed(_zz_10964));
  assign _zz_1505 = _zz_10965[15 : 0];
  assign _zz_2546 = ($signed(_zz_10966) + $signed(_zz_10967));
  assign _zz_1506 = _zz_10968[15 : 0];
  assign _zz_1507 = 1'b1;
  assign _zz_1508 = 1'b1;
  assign _zz_2547 = ($signed(_zz_10985) - $signed(_zz_10986));
  assign _zz_1509 = _zz_10987[15 : 0];
  assign _zz_2548 = ($signed(_zz_10988) + $signed(_zz_10989));
  assign _zz_1510 = _zz_10990[15 : 0];
  assign _zz_1511 = 1'b1;
  assign _zz_1512 = 1'b1;
  assign _zz_2549 = ($signed(_zz_11007) - $signed(_zz_11008));
  assign _zz_1513 = _zz_11009[15 : 0];
  assign _zz_2550 = ($signed(_zz_11010) + $signed(_zz_11011));
  assign _zz_1514 = _zz_11012[15 : 0];
  assign _zz_1515 = 1'b1;
  assign _zz_1516 = 1'b1;
  assign _zz_2551 = ($signed(_zz_11029) - $signed(_zz_11030));
  assign _zz_1517 = _zz_11031[15 : 0];
  assign _zz_2552 = ($signed(_zz_11032) + $signed(_zz_11033));
  assign _zz_1518 = _zz_11034[15 : 0];
  assign _zz_1519 = 1'b1;
  assign _zz_1520 = 1'b1;
  assign _zz_2553 = ($signed(_zz_11051) - $signed(_zz_11052));
  assign _zz_1521 = _zz_11053[15 : 0];
  assign _zz_2554 = ($signed(_zz_11054) + $signed(_zz_11055));
  assign _zz_1522 = _zz_11056[15 : 0];
  assign _zz_1523 = 1'b1;
  assign _zz_1524 = 1'b1;
  assign _zz_2555 = ($signed(_zz_11073) - $signed(_zz_11074));
  assign _zz_1525 = _zz_11075[15 : 0];
  assign _zz_2556 = ($signed(_zz_11076) + $signed(_zz_11077));
  assign _zz_1526 = _zz_11078[15 : 0];
  assign _zz_1527 = 1'b1;
  assign _zz_1528 = 1'b1;
  assign _zz_2557 = ($signed(_zz_11095) - $signed(_zz_11096));
  assign _zz_1529 = _zz_11097[15 : 0];
  assign _zz_2558 = ($signed(_zz_11098) + $signed(_zz_11099));
  assign _zz_1530 = _zz_11100[15 : 0];
  assign _zz_1531 = 1'b1;
  assign _zz_1532 = 1'b1;
  assign _zz_2559 = ($signed(_zz_11117) - $signed(_zz_11118));
  assign _zz_1533 = _zz_11119[15 : 0];
  assign _zz_2560 = ($signed(_zz_11120) + $signed(_zz_11121));
  assign _zz_1534 = _zz_11122[15 : 0];
  assign _zz_1535 = 1'b1;
  assign _zz_1536 = 1'b1;
  assign _zz_2561 = ($signed(_zz_11139) - $signed(_zz_11140));
  assign _zz_1537 = _zz_11141[15 : 0];
  assign _zz_2562 = ($signed(_zz_11142) + $signed(_zz_11143));
  assign _zz_1538 = _zz_11144[15 : 0];
  assign _zz_1539 = 1'b1;
  assign _zz_1540 = 1'b1;
  assign _zz_2563 = ($signed(_zz_11161) - $signed(_zz_11162));
  assign _zz_1541 = _zz_11163[15 : 0];
  assign _zz_2564 = ($signed(_zz_11164) + $signed(_zz_11165));
  assign _zz_1542 = _zz_11166[15 : 0];
  assign _zz_1543 = 1'b1;
  assign _zz_1544 = 1'b1;
  assign _zz_2565 = ($signed(_zz_11183) - $signed(_zz_11184));
  assign _zz_1545 = _zz_11185[15 : 0];
  assign _zz_2566 = ($signed(_zz_11186) + $signed(_zz_11187));
  assign _zz_1546 = _zz_11188[15 : 0];
  assign _zz_1547 = 1'b1;
  assign _zz_1548 = 1'b1;
  assign _zz_2567 = ($signed(_zz_11205) - $signed(_zz_11206));
  assign _zz_1549 = _zz_11207[15 : 0];
  assign _zz_2568 = ($signed(_zz_11208) + $signed(_zz_11209));
  assign _zz_1550 = _zz_11210[15 : 0];
  assign _zz_1551 = 1'b1;
  assign _zz_1552 = 1'b1;
  assign _zz_2569 = ($signed(_zz_11227) - $signed(_zz_11228));
  assign _zz_1553 = _zz_11229[15 : 0];
  assign _zz_2570 = ($signed(_zz_11230) + $signed(_zz_11231));
  assign _zz_1554 = _zz_11232[15 : 0];
  assign _zz_1555 = 1'b1;
  assign _zz_1556 = 1'b1;
  assign _zz_2571 = ($signed(_zz_11249) - $signed(_zz_11250));
  assign _zz_1557 = _zz_11251[15 : 0];
  assign _zz_2572 = ($signed(_zz_11252) + $signed(_zz_11253));
  assign _zz_1558 = _zz_11254[15 : 0];
  assign _zz_1559 = 1'b1;
  assign _zz_1560 = 1'b1;
  assign _zz_2573 = ($signed(_zz_11271) - $signed(_zz_11272));
  assign _zz_1561 = _zz_11273[15 : 0];
  assign _zz_2574 = ($signed(_zz_11274) + $signed(_zz_11275));
  assign _zz_1562 = _zz_11276[15 : 0];
  assign _zz_1563 = 1'b1;
  assign _zz_1564 = 1'b1;
  assign _zz_2575 = ($signed(_zz_11293) - $signed(_zz_11294));
  assign _zz_1565 = _zz_11295[15 : 0];
  assign _zz_2576 = ($signed(_zz_11296) + $signed(_zz_11297));
  assign _zz_1566 = _zz_11298[15 : 0];
  assign _zz_1567 = 1'b1;
  assign _zz_1568 = 1'b1;
  assign _zz_2577 = ($signed(_zz_11315) - $signed(_zz_11316));
  assign _zz_1569 = _zz_11317[15 : 0];
  assign _zz_2578 = ($signed(_zz_11318) + $signed(_zz_11319));
  assign _zz_1570 = _zz_11320[15 : 0];
  assign _zz_1571 = 1'b1;
  assign _zz_1572 = 1'b1;
  assign _zz_2579 = ($signed(_zz_11337) - $signed(_zz_11338));
  assign _zz_1573 = _zz_11339[15 : 0];
  assign _zz_2580 = ($signed(_zz_11340) + $signed(_zz_11341));
  assign _zz_1574 = _zz_11342[15 : 0];
  assign _zz_1575 = 1'b1;
  assign _zz_1576 = 1'b1;
  assign _zz_2581 = ($signed(_zz_11359) - $signed(_zz_11360));
  assign _zz_1577 = _zz_11361[15 : 0];
  assign _zz_2582 = ($signed(_zz_11362) + $signed(_zz_11363));
  assign _zz_1578 = _zz_11364[15 : 0];
  assign _zz_1579 = 1'b1;
  assign _zz_1580 = 1'b1;
  assign _zz_2583 = ($signed(_zz_11381) - $signed(_zz_11382));
  assign _zz_1581 = _zz_11383[15 : 0];
  assign _zz_2584 = ($signed(_zz_11384) + $signed(_zz_11385));
  assign _zz_1582 = _zz_11386[15 : 0];
  assign _zz_1583 = 1'b1;
  assign _zz_1584 = 1'b1;
  assign _zz_2585 = ($signed(_zz_11403) - $signed(_zz_11404));
  assign _zz_1585 = _zz_11405[15 : 0];
  assign _zz_2586 = ($signed(_zz_11406) + $signed(_zz_11407));
  assign _zz_1586 = _zz_11408[15 : 0];
  assign _zz_1587 = 1'b1;
  assign _zz_1588 = 1'b1;
  assign _zz_2587 = ($signed(_zz_11425) - $signed(_zz_11426));
  assign _zz_1589 = _zz_11427[15 : 0];
  assign _zz_2588 = ($signed(_zz_11428) + $signed(_zz_11429));
  assign _zz_1590 = _zz_11430[15 : 0];
  assign _zz_1591 = 1'b1;
  assign _zz_1592 = 1'b1;
  assign _zz_2589 = ($signed(_zz_11447) - $signed(_zz_11448));
  assign _zz_1593 = _zz_11449[15 : 0];
  assign _zz_2590 = ($signed(_zz_11450) + $signed(_zz_11451));
  assign _zz_1594 = _zz_11452[15 : 0];
  assign _zz_1595 = 1'b1;
  assign _zz_1596 = 1'b1;
  assign _zz_2591 = ($signed(_zz_11469) - $signed(_zz_11470));
  assign _zz_1597 = _zz_11471[15 : 0];
  assign _zz_2592 = ($signed(_zz_11472) + $signed(_zz_11473));
  assign _zz_1598 = _zz_11474[15 : 0];
  assign _zz_1599 = 1'b1;
  assign _zz_1600 = 1'b1;
  assign _zz_2593 = ($signed(_zz_11491) - $signed(_zz_11492));
  assign _zz_1601 = _zz_11493[15 : 0];
  assign _zz_2594 = ($signed(_zz_11494) + $signed(_zz_11495));
  assign _zz_1602 = _zz_11496[15 : 0];
  assign _zz_1603 = 1'b1;
  assign _zz_1604 = 1'b1;
  assign _zz_2595 = ($signed(_zz_11513) - $signed(_zz_11514));
  assign _zz_1605 = _zz_11515[15 : 0];
  assign _zz_2596 = ($signed(_zz_11516) + $signed(_zz_11517));
  assign _zz_1606 = _zz_11518[15 : 0];
  assign _zz_1607 = 1'b1;
  assign _zz_1608 = 1'b1;
  assign _zz_2597 = ($signed(_zz_11535) - $signed(_zz_11536));
  assign _zz_1609 = _zz_11537[15 : 0];
  assign _zz_2598 = ($signed(_zz_11538) + $signed(_zz_11539));
  assign _zz_1610 = _zz_11540[15 : 0];
  assign _zz_1611 = 1'b1;
  assign _zz_1612 = 1'b1;
  assign _zz_2599 = ($signed(_zz_11557) - $signed(_zz_11558));
  assign _zz_1613 = _zz_11559[15 : 0];
  assign _zz_2600 = ($signed(_zz_11560) + $signed(_zz_11561));
  assign _zz_1614 = _zz_11562[15 : 0];
  assign _zz_1615 = 1'b1;
  assign _zz_1616 = 1'b1;
  assign _zz_2601 = ($signed(_zz_11579) - $signed(_zz_11580));
  assign _zz_1617 = _zz_11581[15 : 0];
  assign _zz_2602 = ($signed(_zz_11582) + $signed(_zz_11583));
  assign _zz_1618 = _zz_11584[15 : 0];
  assign _zz_1619 = 1'b1;
  assign _zz_1620 = 1'b1;
  assign _zz_2603 = ($signed(_zz_11601) - $signed(_zz_11602));
  assign _zz_1621 = _zz_11603[15 : 0];
  assign _zz_2604 = ($signed(_zz_11604) + $signed(_zz_11605));
  assign _zz_1622 = _zz_11606[15 : 0];
  assign _zz_1623 = 1'b1;
  assign _zz_1624 = 1'b1;
  assign _zz_2605 = ($signed(_zz_11623) - $signed(_zz_11624));
  assign _zz_1625 = _zz_11625[15 : 0];
  assign _zz_2606 = ($signed(_zz_11626) + $signed(_zz_11627));
  assign _zz_1626 = _zz_11628[15 : 0];
  assign _zz_1627 = 1'b1;
  assign _zz_1628 = 1'b1;
  assign _zz_2607 = ($signed(_zz_11645) - $signed(_zz_11646));
  assign _zz_1629 = _zz_11647[15 : 0];
  assign _zz_2608 = ($signed(_zz_11648) + $signed(_zz_11649));
  assign _zz_1630 = _zz_11650[15 : 0];
  assign _zz_1631 = 1'b1;
  assign _zz_1632 = 1'b1;
  assign _zz_2609 = ($signed(_zz_11667) - $signed(_zz_11668));
  assign _zz_1633 = _zz_11669[15 : 0];
  assign _zz_2610 = ($signed(_zz_11670) + $signed(_zz_11671));
  assign _zz_1634 = _zz_11672[15 : 0];
  assign _zz_1635 = 1'b1;
  assign _zz_1636 = 1'b1;
  assign _zz_2611 = ($signed(_zz_11689) - $signed(_zz_11690));
  assign _zz_1637 = _zz_11691[15 : 0];
  assign _zz_2612 = ($signed(_zz_11692) + $signed(_zz_11693));
  assign _zz_1638 = _zz_11694[15 : 0];
  assign _zz_1639 = 1'b1;
  assign _zz_1640 = 1'b1;
  assign _zz_2613 = ($signed(_zz_11711) - $signed(_zz_11712));
  assign _zz_1641 = _zz_11713[15 : 0];
  assign _zz_2614 = ($signed(_zz_11714) + $signed(_zz_11715));
  assign _zz_1642 = _zz_11716[15 : 0];
  assign _zz_1643 = 1'b1;
  assign _zz_1644 = 1'b1;
  assign _zz_2615 = ($signed(_zz_11733) - $signed(_zz_11734));
  assign _zz_1645 = _zz_11735[15 : 0];
  assign _zz_2616 = ($signed(_zz_11736) + $signed(_zz_11737));
  assign _zz_1646 = _zz_11738[15 : 0];
  assign _zz_1647 = 1'b1;
  assign _zz_1648 = 1'b1;
  assign _zz_2617 = ($signed(_zz_11755) - $signed(_zz_11756));
  assign _zz_1649 = _zz_11757[15 : 0];
  assign _zz_2618 = ($signed(_zz_11758) + $signed(_zz_11759));
  assign _zz_1650 = _zz_11760[15 : 0];
  assign _zz_1651 = 1'b1;
  assign _zz_1652 = 1'b1;
  assign _zz_2619 = ($signed(_zz_11777) - $signed(_zz_11778));
  assign _zz_1653 = _zz_11779[15 : 0];
  assign _zz_2620 = ($signed(_zz_11780) + $signed(_zz_11781));
  assign _zz_1654 = _zz_11782[15 : 0];
  assign _zz_1655 = 1'b1;
  assign _zz_1656 = 1'b1;
  assign _zz_2621 = ($signed(_zz_11799) - $signed(_zz_11800));
  assign _zz_1657 = _zz_11801[15 : 0];
  assign _zz_2622 = ($signed(_zz_11802) + $signed(_zz_11803));
  assign _zz_1658 = _zz_11804[15 : 0];
  assign _zz_1659 = 1'b1;
  assign _zz_1660 = 1'b1;
  assign _zz_2623 = ($signed(_zz_11821) - $signed(_zz_11822));
  assign _zz_1661 = _zz_11823[15 : 0];
  assign _zz_2624 = ($signed(_zz_11824) + $signed(_zz_11825));
  assign _zz_1662 = _zz_11826[15 : 0];
  assign _zz_1663 = 1'b1;
  assign _zz_1664 = 1'b1;
  assign _zz_2625 = ($signed(_zz_11843) - $signed(_zz_11844));
  assign _zz_1665 = _zz_11845[15 : 0];
  assign _zz_2626 = ($signed(_zz_11846) + $signed(_zz_11847));
  assign _zz_1666 = _zz_11848[15 : 0];
  assign _zz_1667 = 1'b1;
  assign _zz_1668 = 1'b1;
  assign _zz_2627 = ($signed(_zz_11865) - $signed(_zz_11866));
  assign _zz_1669 = _zz_11867[15 : 0];
  assign _zz_2628 = ($signed(_zz_11868) + $signed(_zz_11869));
  assign _zz_1670 = _zz_11870[15 : 0];
  assign _zz_1671 = 1'b1;
  assign _zz_1672 = 1'b1;
  assign _zz_2629 = ($signed(_zz_11887) - $signed(_zz_11888));
  assign _zz_1673 = _zz_11889[15 : 0];
  assign _zz_2630 = ($signed(_zz_11890) + $signed(_zz_11891));
  assign _zz_1674 = _zz_11892[15 : 0];
  assign _zz_1675 = 1'b1;
  assign _zz_1676 = 1'b1;
  assign _zz_2631 = ($signed(_zz_11909) - $signed(_zz_11910));
  assign _zz_1677 = _zz_11911[15 : 0];
  assign _zz_2632 = ($signed(_zz_11912) + $signed(_zz_11913));
  assign _zz_1678 = _zz_11914[15 : 0];
  assign _zz_1679 = 1'b1;
  assign _zz_1680 = 1'b1;
  assign _zz_2633 = ($signed(_zz_11931) - $signed(_zz_11932));
  assign _zz_1681 = _zz_11933[15 : 0];
  assign _zz_2634 = ($signed(_zz_11934) + $signed(_zz_11935));
  assign _zz_1682 = _zz_11936[15 : 0];
  assign _zz_1683 = 1'b1;
  assign _zz_1684 = 1'b1;
  assign _zz_2635 = ($signed(_zz_11953) - $signed(_zz_11954));
  assign _zz_1685 = _zz_11955[15 : 0];
  assign _zz_2636 = ($signed(_zz_11956) + $signed(_zz_11957));
  assign _zz_1686 = _zz_11958[15 : 0];
  assign _zz_1687 = 1'b1;
  assign _zz_1688 = 1'b1;
  assign _zz_2637 = ($signed(_zz_11975) - $signed(_zz_11976));
  assign _zz_1689 = _zz_11977[15 : 0];
  assign _zz_2638 = ($signed(_zz_11978) + $signed(_zz_11979));
  assign _zz_1690 = _zz_11980[15 : 0];
  assign _zz_1691 = 1'b1;
  assign _zz_1692 = 1'b1;
  assign _zz_2639 = ($signed(_zz_11997) - $signed(_zz_11998));
  assign _zz_1693 = _zz_11999[15 : 0];
  assign _zz_2640 = ($signed(_zz_12000) + $signed(_zz_12001));
  assign _zz_1694 = _zz_12002[15 : 0];
  assign _zz_1695 = 1'b1;
  assign _zz_1696 = 1'b1;
  assign _zz_2641 = ($signed(_zz_12019) - $signed(_zz_12020));
  assign _zz_1697 = _zz_12021[15 : 0];
  assign _zz_2642 = ($signed(_zz_12022) + $signed(_zz_12023));
  assign _zz_1698 = _zz_12024[15 : 0];
  assign _zz_1699 = 1'b1;
  assign _zz_1700 = 1'b1;
  assign _zz_2643 = ($signed(_zz_12041) - $signed(_zz_12042));
  assign _zz_1701 = _zz_12043[15 : 0];
  assign _zz_2644 = ($signed(_zz_12044) + $signed(_zz_12045));
  assign _zz_1702 = _zz_12046[15 : 0];
  assign _zz_1703 = 1'b1;
  assign _zz_1704 = 1'b1;
  assign _zz_2645 = ($signed(_zz_12063) - $signed(_zz_12064));
  assign _zz_1705 = _zz_12065[15 : 0];
  assign _zz_2646 = ($signed(_zz_12066) + $signed(_zz_12067));
  assign _zz_1706 = _zz_12068[15 : 0];
  assign _zz_1707 = 1'b1;
  assign _zz_1708 = 1'b1;
  assign _zz_2647 = ($signed(_zz_12085) - $signed(_zz_12086));
  assign _zz_1709 = _zz_12087[15 : 0];
  assign _zz_2648 = ($signed(_zz_12088) + $signed(_zz_12089));
  assign _zz_1710 = _zz_12090[15 : 0];
  assign _zz_1711 = 1'b1;
  assign _zz_1712 = 1'b1;
  assign _zz_2649 = ($signed(_zz_12107) - $signed(_zz_12108));
  assign _zz_1713 = _zz_12109[15 : 0];
  assign _zz_2650 = ($signed(_zz_12110) + $signed(_zz_12111));
  assign _zz_1714 = _zz_12112[15 : 0];
  assign _zz_1715 = 1'b1;
  assign _zz_1716 = 1'b1;
  assign _zz_2651 = ($signed(_zz_12129) - $signed(_zz_12130));
  assign _zz_1717 = _zz_12131[15 : 0];
  assign _zz_2652 = ($signed(_zz_12132) + $signed(_zz_12133));
  assign _zz_1718 = _zz_12134[15 : 0];
  assign _zz_1719 = 1'b1;
  assign _zz_1720 = 1'b1;
  assign _zz_2653 = ($signed(_zz_12151) - $signed(_zz_12152));
  assign _zz_1721 = _zz_12153[15 : 0];
  assign _zz_2654 = ($signed(_zz_12154) + $signed(_zz_12155));
  assign _zz_1722 = _zz_12156[15 : 0];
  assign _zz_1723 = 1'b1;
  assign _zz_1724 = 1'b1;
  assign _zz_2655 = ($signed(_zz_12173) - $signed(_zz_12174));
  assign _zz_1725 = _zz_12175[15 : 0];
  assign _zz_2656 = ($signed(_zz_12176) + $signed(_zz_12177));
  assign _zz_1726 = _zz_12178[15 : 0];
  assign _zz_1727 = 1'b1;
  assign _zz_1728 = 1'b1;
  assign _zz_2657 = ($signed(_zz_12195) - $signed(_zz_12196));
  assign _zz_1729 = _zz_12197[15 : 0];
  assign _zz_2658 = ($signed(_zz_12198) + $signed(_zz_12199));
  assign _zz_1730 = _zz_12200[15 : 0];
  assign _zz_1731 = 1'b1;
  assign _zz_1732 = 1'b1;
  assign _zz_2659 = ($signed(_zz_12217) - $signed(_zz_12218));
  assign _zz_1733 = _zz_12219[15 : 0];
  assign _zz_2660 = ($signed(_zz_12220) + $signed(_zz_12221));
  assign _zz_1734 = _zz_12222[15 : 0];
  assign _zz_1735 = 1'b1;
  assign _zz_1736 = 1'b1;
  assign _zz_2661 = ($signed(_zz_12239) - $signed(_zz_12240));
  assign _zz_1737 = _zz_12241[15 : 0];
  assign _zz_2662 = ($signed(_zz_12242) + $signed(_zz_12243));
  assign _zz_1738 = _zz_12244[15 : 0];
  assign _zz_1739 = 1'b1;
  assign _zz_1740 = 1'b1;
  assign _zz_2663 = ($signed(_zz_12261) - $signed(_zz_12262));
  assign _zz_1741 = _zz_12263[15 : 0];
  assign _zz_2664 = ($signed(_zz_12264) + $signed(_zz_12265));
  assign _zz_1742 = _zz_12266[15 : 0];
  assign _zz_1743 = 1'b1;
  assign _zz_1744 = 1'b1;
  assign _zz_2665 = ($signed(_zz_12283) - $signed(_zz_12284));
  assign _zz_1745 = _zz_12285[15 : 0];
  assign _zz_2666 = ($signed(_zz_12286) + $signed(_zz_12287));
  assign _zz_1746 = _zz_12288[15 : 0];
  assign _zz_1747 = 1'b1;
  assign _zz_1748 = 1'b1;
  assign _zz_2667 = ($signed(_zz_12305) - $signed(_zz_12306));
  assign _zz_1749 = _zz_12307[15 : 0];
  assign _zz_2668 = ($signed(_zz_12308) + $signed(_zz_12309));
  assign _zz_1750 = _zz_12310[15 : 0];
  assign _zz_1751 = 1'b1;
  assign _zz_1752 = 1'b1;
  assign _zz_2669 = ($signed(_zz_12327) - $signed(_zz_12328));
  assign _zz_1753 = _zz_12329[15 : 0];
  assign _zz_2670 = ($signed(_zz_12330) + $signed(_zz_12331));
  assign _zz_1754 = _zz_12332[15 : 0];
  assign _zz_1755 = 1'b1;
  assign _zz_1756 = 1'b1;
  assign _zz_2671 = ($signed(_zz_12349) - $signed(_zz_12350));
  assign _zz_1757 = _zz_12351[15 : 0];
  assign _zz_2672 = ($signed(_zz_12352) + $signed(_zz_12353));
  assign _zz_1758 = _zz_12354[15 : 0];
  assign _zz_1759 = 1'b1;
  assign _zz_1760 = 1'b1;
  assign _zz_2673 = ($signed(_zz_12371) - $signed(_zz_12372));
  assign _zz_1761 = _zz_12373[15 : 0];
  assign _zz_2674 = ($signed(_zz_12374) + $signed(_zz_12375));
  assign _zz_1762 = _zz_12376[15 : 0];
  assign _zz_1763 = 1'b1;
  assign _zz_1764 = 1'b1;
  assign _zz_2675 = ($signed(_zz_12393) - $signed(_zz_12394));
  assign _zz_1765 = _zz_12395[15 : 0];
  assign _zz_2676 = ($signed(_zz_12396) + $signed(_zz_12397));
  assign _zz_1766 = _zz_12398[15 : 0];
  assign _zz_1767 = 1'b1;
  assign _zz_1768 = 1'b1;
  assign _zz_2677 = ($signed(_zz_12415) - $signed(_zz_12416));
  assign _zz_1769 = _zz_12417[15 : 0];
  assign _zz_2678 = ($signed(_zz_12418) + $signed(_zz_12419));
  assign _zz_1770 = _zz_12420[15 : 0];
  assign _zz_1771 = 1'b1;
  assign _zz_1772 = 1'b1;
  assign _zz_2679 = ($signed(_zz_12437) - $signed(_zz_12438));
  assign _zz_1773 = _zz_12439[15 : 0];
  assign _zz_2680 = ($signed(_zz_12440) + $signed(_zz_12441));
  assign _zz_1774 = _zz_12442[15 : 0];
  assign _zz_1775 = 1'b1;
  assign _zz_1776 = 1'b1;
  assign _zz_2681 = ($signed(_zz_12459) - $signed(_zz_12460));
  assign _zz_1777 = _zz_12461[15 : 0];
  assign _zz_2682 = ($signed(_zz_12462) + $signed(_zz_12463));
  assign _zz_1778 = _zz_12464[15 : 0];
  assign _zz_1779 = 1'b1;
  assign _zz_1780 = 1'b1;
  assign _zz_2683 = ($signed(_zz_12481) - $signed(_zz_12482));
  assign _zz_1781 = _zz_12483[15 : 0];
  assign _zz_2684 = ($signed(_zz_12484) + $signed(_zz_12485));
  assign _zz_1782 = _zz_12486[15 : 0];
  assign _zz_1783 = 1'b1;
  assign _zz_1784 = 1'b1;
  assign _zz_2685 = ($signed(_zz_12503) - $signed(_zz_12504));
  assign _zz_1785 = _zz_12505[15 : 0];
  assign _zz_2686 = ($signed(_zz_12506) + $signed(_zz_12507));
  assign _zz_1786 = _zz_12508[15 : 0];
  assign _zz_1787 = 1'b1;
  assign _zz_1788 = 1'b1;
  assign _zz_2687 = ($signed(_zz_12525) - $signed(_zz_12526));
  assign _zz_1789 = _zz_12527[15 : 0];
  assign _zz_2688 = ($signed(_zz_12528) + $signed(_zz_12529));
  assign _zz_1790 = _zz_12530[15 : 0];
  assign _zz_1791 = 1'b1;
  assign _zz_1792 = 1'b1;
  assign io_data_out_valid = current_level_cnt_willOverflow_regNext;
  assign io_data_out_payload_0_real = data_mid_0_real;
  assign io_data_out_payload_0_imag = data_mid_0_imag;
  assign io_data_out_payload_1_real = data_mid_1_real;
  assign io_data_out_payload_1_imag = data_mid_1_imag;
  assign io_data_out_payload_2_real = data_mid_2_real;
  assign io_data_out_payload_2_imag = data_mid_2_imag;
  assign io_data_out_payload_3_real = data_mid_3_real;
  assign io_data_out_payload_3_imag = data_mid_3_imag;
  assign io_data_out_payload_4_real = data_mid_4_real;
  assign io_data_out_payload_4_imag = data_mid_4_imag;
  assign io_data_out_payload_5_real = data_mid_5_real;
  assign io_data_out_payload_5_imag = data_mid_5_imag;
  assign io_data_out_payload_6_real = data_mid_6_real;
  assign io_data_out_payload_6_imag = data_mid_6_imag;
  assign io_data_out_payload_7_real = data_mid_7_real;
  assign io_data_out_payload_7_imag = data_mid_7_imag;
  assign io_data_out_payload_8_real = data_mid_8_real;
  assign io_data_out_payload_8_imag = data_mid_8_imag;
  assign io_data_out_payload_9_real = data_mid_9_real;
  assign io_data_out_payload_9_imag = data_mid_9_imag;
  assign io_data_out_payload_10_real = data_mid_10_real;
  assign io_data_out_payload_10_imag = data_mid_10_imag;
  assign io_data_out_payload_11_real = data_mid_11_real;
  assign io_data_out_payload_11_imag = data_mid_11_imag;
  assign io_data_out_payload_12_real = data_mid_12_real;
  assign io_data_out_payload_12_imag = data_mid_12_imag;
  assign io_data_out_payload_13_real = data_mid_13_real;
  assign io_data_out_payload_13_imag = data_mid_13_imag;
  assign io_data_out_payload_14_real = data_mid_14_real;
  assign io_data_out_payload_14_imag = data_mid_14_imag;
  assign io_data_out_payload_15_real = data_mid_15_real;
  assign io_data_out_payload_15_imag = data_mid_15_imag;
  assign io_data_out_payload_16_real = data_mid_16_real;
  assign io_data_out_payload_16_imag = data_mid_16_imag;
  assign io_data_out_payload_17_real = data_mid_17_real;
  assign io_data_out_payload_17_imag = data_mid_17_imag;
  assign io_data_out_payload_18_real = data_mid_18_real;
  assign io_data_out_payload_18_imag = data_mid_18_imag;
  assign io_data_out_payload_19_real = data_mid_19_real;
  assign io_data_out_payload_19_imag = data_mid_19_imag;
  assign io_data_out_payload_20_real = data_mid_20_real;
  assign io_data_out_payload_20_imag = data_mid_20_imag;
  assign io_data_out_payload_21_real = data_mid_21_real;
  assign io_data_out_payload_21_imag = data_mid_21_imag;
  assign io_data_out_payload_22_real = data_mid_22_real;
  assign io_data_out_payload_22_imag = data_mid_22_imag;
  assign io_data_out_payload_23_real = data_mid_23_real;
  assign io_data_out_payload_23_imag = data_mid_23_imag;
  assign io_data_out_payload_24_real = data_mid_24_real;
  assign io_data_out_payload_24_imag = data_mid_24_imag;
  assign io_data_out_payload_25_real = data_mid_25_real;
  assign io_data_out_payload_25_imag = data_mid_25_imag;
  assign io_data_out_payload_26_real = data_mid_26_real;
  assign io_data_out_payload_26_imag = data_mid_26_imag;
  assign io_data_out_payload_27_real = data_mid_27_real;
  assign io_data_out_payload_27_imag = data_mid_27_imag;
  assign io_data_out_payload_28_real = data_mid_28_real;
  assign io_data_out_payload_28_imag = data_mid_28_imag;
  assign io_data_out_payload_29_real = data_mid_29_real;
  assign io_data_out_payload_29_imag = data_mid_29_imag;
  assign io_data_out_payload_30_real = data_mid_30_real;
  assign io_data_out_payload_30_imag = data_mid_30_imag;
  assign io_data_out_payload_31_real = data_mid_31_real;
  assign io_data_out_payload_31_imag = data_mid_31_imag;
  assign io_data_out_payload_32_real = data_mid_32_real;
  assign io_data_out_payload_32_imag = data_mid_32_imag;
  assign io_data_out_payload_33_real = data_mid_33_real;
  assign io_data_out_payload_33_imag = data_mid_33_imag;
  assign io_data_out_payload_34_real = data_mid_34_real;
  assign io_data_out_payload_34_imag = data_mid_34_imag;
  assign io_data_out_payload_35_real = data_mid_35_real;
  assign io_data_out_payload_35_imag = data_mid_35_imag;
  assign io_data_out_payload_36_real = data_mid_36_real;
  assign io_data_out_payload_36_imag = data_mid_36_imag;
  assign io_data_out_payload_37_real = data_mid_37_real;
  assign io_data_out_payload_37_imag = data_mid_37_imag;
  assign io_data_out_payload_38_real = data_mid_38_real;
  assign io_data_out_payload_38_imag = data_mid_38_imag;
  assign io_data_out_payload_39_real = data_mid_39_real;
  assign io_data_out_payload_39_imag = data_mid_39_imag;
  assign io_data_out_payload_40_real = data_mid_40_real;
  assign io_data_out_payload_40_imag = data_mid_40_imag;
  assign io_data_out_payload_41_real = data_mid_41_real;
  assign io_data_out_payload_41_imag = data_mid_41_imag;
  assign io_data_out_payload_42_real = data_mid_42_real;
  assign io_data_out_payload_42_imag = data_mid_42_imag;
  assign io_data_out_payload_43_real = data_mid_43_real;
  assign io_data_out_payload_43_imag = data_mid_43_imag;
  assign io_data_out_payload_44_real = data_mid_44_real;
  assign io_data_out_payload_44_imag = data_mid_44_imag;
  assign io_data_out_payload_45_real = data_mid_45_real;
  assign io_data_out_payload_45_imag = data_mid_45_imag;
  assign io_data_out_payload_46_real = data_mid_46_real;
  assign io_data_out_payload_46_imag = data_mid_46_imag;
  assign io_data_out_payload_47_real = data_mid_47_real;
  assign io_data_out_payload_47_imag = data_mid_47_imag;
  assign io_data_out_payload_48_real = data_mid_48_real;
  assign io_data_out_payload_48_imag = data_mid_48_imag;
  assign io_data_out_payload_49_real = data_mid_49_real;
  assign io_data_out_payload_49_imag = data_mid_49_imag;
  assign io_data_out_payload_50_real = data_mid_50_real;
  assign io_data_out_payload_50_imag = data_mid_50_imag;
  assign io_data_out_payload_51_real = data_mid_51_real;
  assign io_data_out_payload_51_imag = data_mid_51_imag;
  assign io_data_out_payload_52_real = data_mid_52_real;
  assign io_data_out_payload_52_imag = data_mid_52_imag;
  assign io_data_out_payload_53_real = data_mid_53_real;
  assign io_data_out_payload_53_imag = data_mid_53_imag;
  assign io_data_out_payload_54_real = data_mid_54_real;
  assign io_data_out_payload_54_imag = data_mid_54_imag;
  assign io_data_out_payload_55_real = data_mid_55_real;
  assign io_data_out_payload_55_imag = data_mid_55_imag;
  assign io_data_out_payload_56_real = data_mid_56_real;
  assign io_data_out_payload_56_imag = data_mid_56_imag;
  assign io_data_out_payload_57_real = data_mid_57_real;
  assign io_data_out_payload_57_imag = data_mid_57_imag;
  assign io_data_out_payload_58_real = data_mid_58_real;
  assign io_data_out_payload_58_imag = data_mid_58_imag;
  assign io_data_out_payload_59_real = data_mid_59_real;
  assign io_data_out_payload_59_imag = data_mid_59_imag;
  assign io_data_out_payload_60_real = data_mid_60_real;
  assign io_data_out_payload_60_imag = data_mid_60_imag;
  assign io_data_out_payload_61_real = data_mid_61_real;
  assign io_data_out_payload_61_imag = data_mid_61_imag;
  assign io_data_out_payload_62_real = data_mid_62_real;
  assign io_data_out_payload_62_imag = data_mid_62_imag;
  assign io_data_out_payload_63_real = data_mid_63_real;
  assign io_data_out_payload_63_imag = data_mid_63_imag;
  assign io_data_out_payload_64_real = data_mid_64_real;
  assign io_data_out_payload_64_imag = data_mid_64_imag;
  assign io_data_out_payload_65_real = data_mid_65_real;
  assign io_data_out_payload_65_imag = data_mid_65_imag;
  assign io_data_out_payload_66_real = data_mid_66_real;
  assign io_data_out_payload_66_imag = data_mid_66_imag;
  assign io_data_out_payload_67_real = data_mid_67_real;
  assign io_data_out_payload_67_imag = data_mid_67_imag;
  assign io_data_out_payload_68_real = data_mid_68_real;
  assign io_data_out_payload_68_imag = data_mid_68_imag;
  assign io_data_out_payload_69_real = data_mid_69_real;
  assign io_data_out_payload_69_imag = data_mid_69_imag;
  assign io_data_out_payload_70_real = data_mid_70_real;
  assign io_data_out_payload_70_imag = data_mid_70_imag;
  assign io_data_out_payload_71_real = data_mid_71_real;
  assign io_data_out_payload_71_imag = data_mid_71_imag;
  assign io_data_out_payload_72_real = data_mid_72_real;
  assign io_data_out_payload_72_imag = data_mid_72_imag;
  assign io_data_out_payload_73_real = data_mid_73_real;
  assign io_data_out_payload_73_imag = data_mid_73_imag;
  assign io_data_out_payload_74_real = data_mid_74_real;
  assign io_data_out_payload_74_imag = data_mid_74_imag;
  assign io_data_out_payload_75_real = data_mid_75_real;
  assign io_data_out_payload_75_imag = data_mid_75_imag;
  assign io_data_out_payload_76_real = data_mid_76_real;
  assign io_data_out_payload_76_imag = data_mid_76_imag;
  assign io_data_out_payload_77_real = data_mid_77_real;
  assign io_data_out_payload_77_imag = data_mid_77_imag;
  assign io_data_out_payload_78_real = data_mid_78_real;
  assign io_data_out_payload_78_imag = data_mid_78_imag;
  assign io_data_out_payload_79_real = data_mid_79_real;
  assign io_data_out_payload_79_imag = data_mid_79_imag;
  assign io_data_out_payload_80_real = data_mid_80_real;
  assign io_data_out_payload_80_imag = data_mid_80_imag;
  assign io_data_out_payload_81_real = data_mid_81_real;
  assign io_data_out_payload_81_imag = data_mid_81_imag;
  assign io_data_out_payload_82_real = data_mid_82_real;
  assign io_data_out_payload_82_imag = data_mid_82_imag;
  assign io_data_out_payload_83_real = data_mid_83_real;
  assign io_data_out_payload_83_imag = data_mid_83_imag;
  assign io_data_out_payload_84_real = data_mid_84_real;
  assign io_data_out_payload_84_imag = data_mid_84_imag;
  assign io_data_out_payload_85_real = data_mid_85_real;
  assign io_data_out_payload_85_imag = data_mid_85_imag;
  assign io_data_out_payload_86_real = data_mid_86_real;
  assign io_data_out_payload_86_imag = data_mid_86_imag;
  assign io_data_out_payload_87_real = data_mid_87_real;
  assign io_data_out_payload_87_imag = data_mid_87_imag;
  assign io_data_out_payload_88_real = data_mid_88_real;
  assign io_data_out_payload_88_imag = data_mid_88_imag;
  assign io_data_out_payload_89_real = data_mid_89_real;
  assign io_data_out_payload_89_imag = data_mid_89_imag;
  assign io_data_out_payload_90_real = data_mid_90_real;
  assign io_data_out_payload_90_imag = data_mid_90_imag;
  assign io_data_out_payload_91_real = data_mid_91_real;
  assign io_data_out_payload_91_imag = data_mid_91_imag;
  assign io_data_out_payload_92_real = data_mid_92_real;
  assign io_data_out_payload_92_imag = data_mid_92_imag;
  assign io_data_out_payload_93_real = data_mid_93_real;
  assign io_data_out_payload_93_imag = data_mid_93_imag;
  assign io_data_out_payload_94_real = data_mid_94_real;
  assign io_data_out_payload_94_imag = data_mid_94_imag;
  assign io_data_out_payload_95_real = data_mid_95_real;
  assign io_data_out_payload_95_imag = data_mid_95_imag;
  assign io_data_out_payload_96_real = data_mid_96_real;
  assign io_data_out_payload_96_imag = data_mid_96_imag;
  assign io_data_out_payload_97_real = data_mid_97_real;
  assign io_data_out_payload_97_imag = data_mid_97_imag;
  assign io_data_out_payload_98_real = data_mid_98_real;
  assign io_data_out_payload_98_imag = data_mid_98_imag;
  assign io_data_out_payload_99_real = data_mid_99_real;
  assign io_data_out_payload_99_imag = data_mid_99_imag;
  assign io_data_out_payload_100_real = data_mid_100_real;
  assign io_data_out_payload_100_imag = data_mid_100_imag;
  assign io_data_out_payload_101_real = data_mid_101_real;
  assign io_data_out_payload_101_imag = data_mid_101_imag;
  assign io_data_out_payload_102_real = data_mid_102_real;
  assign io_data_out_payload_102_imag = data_mid_102_imag;
  assign io_data_out_payload_103_real = data_mid_103_real;
  assign io_data_out_payload_103_imag = data_mid_103_imag;
  assign io_data_out_payload_104_real = data_mid_104_real;
  assign io_data_out_payload_104_imag = data_mid_104_imag;
  assign io_data_out_payload_105_real = data_mid_105_real;
  assign io_data_out_payload_105_imag = data_mid_105_imag;
  assign io_data_out_payload_106_real = data_mid_106_real;
  assign io_data_out_payload_106_imag = data_mid_106_imag;
  assign io_data_out_payload_107_real = data_mid_107_real;
  assign io_data_out_payload_107_imag = data_mid_107_imag;
  assign io_data_out_payload_108_real = data_mid_108_real;
  assign io_data_out_payload_108_imag = data_mid_108_imag;
  assign io_data_out_payload_109_real = data_mid_109_real;
  assign io_data_out_payload_109_imag = data_mid_109_imag;
  assign io_data_out_payload_110_real = data_mid_110_real;
  assign io_data_out_payload_110_imag = data_mid_110_imag;
  assign io_data_out_payload_111_real = data_mid_111_real;
  assign io_data_out_payload_111_imag = data_mid_111_imag;
  assign io_data_out_payload_112_real = data_mid_112_real;
  assign io_data_out_payload_112_imag = data_mid_112_imag;
  assign io_data_out_payload_113_real = data_mid_113_real;
  assign io_data_out_payload_113_imag = data_mid_113_imag;
  assign io_data_out_payload_114_real = data_mid_114_real;
  assign io_data_out_payload_114_imag = data_mid_114_imag;
  assign io_data_out_payload_115_real = data_mid_115_real;
  assign io_data_out_payload_115_imag = data_mid_115_imag;
  assign io_data_out_payload_116_real = data_mid_116_real;
  assign io_data_out_payload_116_imag = data_mid_116_imag;
  assign io_data_out_payload_117_real = data_mid_117_real;
  assign io_data_out_payload_117_imag = data_mid_117_imag;
  assign io_data_out_payload_118_real = data_mid_118_real;
  assign io_data_out_payload_118_imag = data_mid_118_imag;
  assign io_data_out_payload_119_real = data_mid_119_real;
  assign io_data_out_payload_119_imag = data_mid_119_imag;
  assign io_data_out_payload_120_real = data_mid_120_real;
  assign io_data_out_payload_120_imag = data_mid_120_imag;
  assign io_data_out_payload_121_real = data_mid_121_real;
  assign io_data_out_payload_121_imag = data_mid_121_imag;
  assign io_data_out_payload_122_real = data_mid_122_real;
  assign io_data_out_payload_122_imag = data_mid_122_imag;
  assign io_data_out_payload_123_real = data_mid_123_real;
  assign io_data_out_payload_123_imag = data_mid_123_imag;
  assign io_data_out_payload_124_real = data_mid_124_real;
  assign io_data_out_payload_124_imag = data_mid_124_imag;
  assign io_data_out_payload_125_real = data_mid_125_real;
  assign io_data_out_payload_125_imag = data_mid_125_imag;
  assign io_data_out_payload_126_real = data_mid_126_real;
  assign io_data_out_payload_126_imag = data_mid_126_imag;
  assign io_data_out_payload_127_real = data_mid_127_real;
  assign io_data_out_payload_127_imag = data_mid_127_imag;
  always @ (posedge clk) begin
    if(io_data_in_valid)begin
      data_in_0_real <= io_data_in_payload_0_real;
      data_in_0_imag <= io_data_in_payload_0_imag;
      data_in_1_real <= io_data_in_payload_1_real;
      data_in_1_imag <= io_data_in_payload_1_imag;
      data_in_2_real <= io_data_in_payload_2_real;
      data_in_2_imag <= io_data_in_payload_2_imag;
      data_in_3_real <= io_data_in_payload_3_real;
      data_in_3_imag <= io_data_in_payload_3_imag;
      data_in_4_real <= io_data_in_payload_4_real;
      data_in_4_imag <= io_data_in_payload_4_imag;
      data_in_5_real <= io_data_in_payload_5_real;
      data_in_5_imag <= io_data_in_payload_5_imag;
      data_in_6_real <= io_data_in_payload_6_real;
      data_in_6_imag <= io_data_in_payload_6_imag;
      data_in_7_real <= io_data_in_payload_7_real;
      data_in_7_imag <= io_data_in_payload_7_imag;
      data_in_8_real <= io_data_in_payload_8_real;
      data_in_8_imag <= io_data_in_payload_8_imag;
      data_in_9_real <= io_data_in_payload_9_real;
      data_in_9_imag <= io_data_in_payload_9_imag;
      data_in_10_real <= io_data_in_payload_10_real;
      data_in_10_imag <= io_data_in_payload_10_imag;
      data_in_11_real <= io_data_in_payload_11_real;
      data_in_11_imag <= io_data_in_payload_11_imag;
      data_in_12_real <= io_data_in_payload_12_real;
      data_in_12_imag <= io_data_in_payload_12_imag;
      data_in_13_real <= io_data_in_payload_13_real;
      data_in_13_imag <= io_data_in_payload_13_imag;
      data_in_14_real <= io_data_in_payload_14_real;
      data_in_14_imag <= io_data_in_payload_14_imag;
      data_in_15_real <= io_data_in_payload_15_real;
      data_in_15_imag <= io_data_in_payload_15_imag;
      data_in_16_real <= io_data_in_payload_16_real;
      data_in_16_imag <= io_data_in_payload_16_imag;
      data_in_17_real <= io_data_in_payload_17_real;
      data_in_17_imag <= io_data_in_payload_17_imag;
      data_in_18_real <= io_data_in_payload_18_real;
      data_in_18_imag <= io_data_in_payload_18_imag;
      data_in_19_real <= io_data_in_payload_19_real;
      data_in_19_imag <= io_data_in_payload_19_imag;
      data_in_20_real <= io_data_in_payload_20_real;
      data_in_20_imag <= io_data_in_payload_20_imag;
      data_in_21_real <= io_data_in_payload_21_real;
      data_in_21_imag <= io_data_in_payload_21_imag;
      data_in_22_real <= io_data_in_payload_22_real;
      data_in_22_imag <= io_data_in_payload_22_imag;
      data_in_23_real <= io_data_in_payload_23_real;
      data_in_23_imag <= io_data_in_payload_23_imag;
      data_in_24_real <= io_data_in_payload_24_real;
      data_in_24_imag <= io_data_in_payload_24_imag;
      data_in_25_real <= io_data_in_payload_25_real;
      data_in_25_imag <= io_data_in_payload_25_imag;
      data_in_26_real <= io_data_in_payload_26_real;
      data_in_26_imag <= io_data_in_payload_26_imag;
      data_in_27_real <= io_data_in_payload_27_real;
      data_in_27_imag <= io_data_in_payload_27_imag;
      data_in_28_real <= io_data_in_payload_28_real;
      data_in_28_imag <= io_data_in_payload_28_imag;
      data_in_29_real <= io_data_in_payload_29_real;
      data_in_29_imag <= io_data_in_payload_29_imag;
      data_in_30_real <= io_data_in_payload_30_real;
      data_in_30_imag <= io_data_in_payload_30_imag;
      data_in_31_real <= io_data_in_payload_31_real;
      data_in_31_imag <= io_data_in_payload_31_imag;
      data_in_32_real <= io_data_in_payload_32_real;
      data_in_32_imag <= io_data_in_payload_32_imag;
      data_in_33_real <= io_data_in_payload_33_real;
      data_in_33_imag <= io_data_in_payload_33_imag;
      data_in_34_real <= io_data_in_payload_34_real;
      data_in_34_imag <= io_data_in_payload_34_imag;
      data_in_35_real <= io_data_in_payload_35_real;
      data_in_35_imag <= io_data_in_payload_35_imag;
      data_in_36_real <= io_data_in_payload_36_real;
      data_in_36_imag <= io_data_in_payload_36_imag;
      data_in_37_real <= io_data_in_payload_37_real;
      data_in_37_imag <= io_data_in_payload_37_imag;
      data_in_38_real <= io_data_in_payload_38_real;
      data_in_38_imag <= io_data_in_payload_38_imag;
      data_in_39_real <= io_data_in_payload_39_real;
      data_in_39_imag <= io_data_in_payload_39_imag;
      data_in_40_real <= io_data_in_payload_40_real;
      data_in_40_imag <= io_data_in_payload_40_imag;
      data_in_41_real <= io_data_in_payload_41_real;
      data_in_41_imag <= io_data_in_payload_41_imag;
      data_in_42_real <= io_data_in_payload_42_real;
      data_in_42_imag <= io_data_in_payload_42_imag;
      data_in_43_real <= io_data_in_payload_43_real;
      data_in_43_imag <= io_data_in_payload_43_imag;
      data_in_44_real <= io_data_in_payload_44_real;
      data_in_44_imag <= io_data_in_payload_44_imag;
      data_in_45_real <= io_data_in_payload_45_real;
      data_in_45_imag <= io_data_in_payload_45_imag;
      data_in_46_real <= io_data_in_payload_46_real;
      data_in_46_imag <= io_data_in_payload_46_imag;
      data_in_47_real <= io_data_in_payload_47_real;
      data_in_47_imag <= io_data_in_payload_47_imag;
      data_in_48_real <= io_data_in_payload_48_real;
      data_in_48_imag <= io_data_in_payload_48_imag;
      data_in_49_real <= io_data_in_payload_49_real;
      data_in_49_imag <= io_data_in_payload_49_imag;
      data_in_50_real <= io_data_in_payload_50_real;
      data_in_50_imag <= io_data_in_payload_50_imag;
      data_in_51_real <= io_data_in_payload_51_real;
      data_in_51_imag <= io_data_in_payload_51_imag;
      data_in_52_real <= io_data_in_payload_52_real;
      data_in_52_imag <= io_data_in_payload_52_imag;
      data_in_53_real <= io_data_in_payload_53_real;
      data_in_53_imag <= io_data_in_payload_53_imag;
      data_in_54_real <= io_data_in_payload_54_real;
      data_in_54_imag <= io_data_in_payload_54_imag;
      data_in_55_real <= io_data_in_payload_55_real;
      data_in_55_imag <= io_data_in_payload_55_imag;
      data_in_56_real <= io_data_in_payload_56_real;
      data_in_56_imag <= io_data_in_payload_56_imag;
      data_in_57_real <= io_data_in_payload_57_real;
      data_in_57_imag <= io_data_in_payload_57_imag;
      data_in_58_real <= io_data_in_payload_58_real;
      data_in_58_imag <= io_data_in_payload_58_imag;
      data_in_59_real <= io_data_in_payload_59_real;
      data_in_59_imag <= io_data_in_payload_59_imag;
      data_in_60_real <= io_data_in_payload_60_real;
      data_in_60_imag <= io_data_in_payload_60_imag;
      data_in_61_real <= io_data_in_payload_61_real;
      data_in_61_imag <= io_data_in_payload_61_imag;
      data_in_62_real <= io_data_in_payload_62_real;
      data_in_62_imag <= io_data_in_payload_62_imag;
      data_in_63_real <= io_data_in_payload_63_real;
      data_in_63_imag <= io_data_in_payload_63_imag;
      data_in_64_real <= io_data_in_payload_64_real;
      data_in_64_imag <= io_data_in_payload_64_imag;
      data_in_65_real <= io_data_in_payload_65_real;
      data_in_65_imag <= io_data_in_payload_65_imag;
      data_in_66_real <= io_data_in_payload_66_real;
      data_in_66_imag <= io_data_in_payload_66_imag;
      data_in_67_real <= io_data_in_payload_67_real;
      data_in_67_imag <= io_data_in_payload_67_imag;
      data_in_68_real <= io_data_in_payload_68_real;
      data_in_68_imag <= io_data_in_payload_68_imag;
      data_in_69_real <= io_data_in_payload_69_real;
      data_in_69_imag <= io_data_in_payload_69_imag;
      data_in_70_real <= io_data_in_payload_70_real;
      data_in_70_imag <= io_data_in_payload_70_imag;
      data_in_71_real <= io_data_in_payload_71_real;
      data_in_71_imag <= io_data_in_payload_71_imag;
      data_in_72_real <= io_data_in_payload_72_real;
      data_in_72_imag <= io_data_in_payload_72_imag;
      data_in_73_real <= io_data_in_payload_73_real;
      data_in_73_imag <= io_data_in_payload_73_imag;
      data_in_74_real <= io_data_in_payload_74_real;
      data_in_74_imag <= io_data_in_payload_74_imag;
      data_in_75_real <= io_data_in_payload_75_real;
      data_in_75_imag <= io_data_in_payload_75_imag;
      data_in_76_real <= io_data_in_payload_76_real;
      data_in_76_imag <= io_data_in_payload_76_imag;
      data_in_77_real <= io_data_in_payload_77_real;
      data_in_77_imag <= io_data_in_payload_77_imag;
      data_in_78_real <= io_data_in_payload_78_real;
      data_in_78_imag <= io_data_in_payload_78_imag;
      data_in_79_real <= io_data_in_payload_79_real;
      data_in_79_imag <= io_data_in_payload_79_imag;
      data_in_80_real <= io_data_in_payload_80_real;
      data_in_80_imag <= io_data_in_payload_80_imag;
      data_in_81_real <= io_data_in_payload_81_real;
      data_in_81_imag <= io_data_in_payload_81_imag;
      data_in_82_real <= io_data_in_payload_82_real;
      data_in_82_imag <= io_data_in_payload_82_imag;
      data_in_83_real <= io_data_in_payload_83_real;
      data_in_83_imag <= io_data_in_payload_83_imag;
      data_in_84_real <= io_data_in_payload_84_real;
      data_in_84_imag <= io_data_in_payload_84_imag;
      data_in_85_real <= io_data_in_payload_85_real;
      data_in_85_imag <= io_data_in_payload_85_imag;
      data_in_86_real <= io_data_in_payload_86_real;
      data_in_86_imag <= io_data_in_payload_86_imag;
      data_in_87_real <= io_data_in_payload_87_real;
      data_in_87_imag <= io_data_in_payload_87_imag;
      data_in_88_real <= io_data_in_payload_88_real;
      data_in_88_imag <= io_data_in_payload_88_imag;
      data_in_89_real <= io_data_in_payload_89_real;
      data_in_89_imag <= io_data_in_payload_89_imag;
      data_in_90_real <= io_data_in_payload_90_real;
      data_in_90_imag <= io_data_in_payload_90_imag;
      data_in_91_real <= io_data_in_payload_91_real;
      data_in_91_imag <= io_data_in_payload_91_imag;
      data_in_92_real <= io_data_in_payload_92_real;
      data_in_92_imag <= io_data_in_payload_92_imag;
      data_in_93_real <= io_data_in_payload_93_real;
      data_in_93_imag <= io_data_in_payload_93_imag;
      data_in_94_real <= io_data_in_payload_94_real;
      data_in_94_imag <= io_data_in_payload_94_imag;
      data_in_95_real <= io_data_in_payload_95_real;
      data_in_95_imag <= io_data_in_payload_95_imag;
      data_in_96_real <= io_data_in_payload_96_real;
      data_in_96_imag <= io_data_in_payload_96_imag;
      data_in_97_real <= io_data_in_payload_97_real;
      data_in_97_imag <= io_data_in_payload_97_imag;
      data_in_98_real <= io_data_in_payload_98_real;
      data_in_98_imag <= io_data_in_payload_98_imag;
      data_in_99_real <= io_data_in_payload_99_real;
      data_in_99_imag <= io_data_in_payload_99_imag;
      data_in_100_real <= io_data_in_payload_100_real;
      data_in_100_imag <= io_data_in_payload_100_imag;
      data_in_101_real <= io_data_in_payload_101_real;
      data_in_101_imag <= io_data_in_payload_101_imag;
      data_in_102_real <= io_data_in_payload_102_real;
      data_in_102_imag <= io_data_in_payload_102_imag;
      data_in_103_real <= io_data_in_payload_103_real;
      data_in_103_imag <= io_data_in_payload_103_imag;
      data_in_104_real <= io_data_in_payload_104_real;
      data_in_104_imag <= io_data_in_payload_104_imag;
      data_in_105_real <= io_data_in_payload_105_real;
      data_in_105_imag <= io_data_in_payload_105_imag;
      data_in_106_real <= io_data_in_payload_106_real;
      data_in_106_imag <= io_data_in_payload_106_imag;
      data_in_107_real <= io_data_in_payload_107_real;
      data_in_107_imag <= io_data_in_payload_107_imag;
      data_in_108_real <= io_data_in_payload_108_real;
      data_in_108_imag <= io_data_in_payload_108_imag;
      data_in_109_real <= io_data_in_payload_109_real;
      data_in_109_imag <= io_data_in_payload_109_imag;
      data_in_110_real <= io_data_in_payload_110_real;
      data_in_110_imag <= io_data_in_payload_110_imag;
      data_in_111_real <= io_data_in_payload_111_real;
      data_in_111_imag <= io_data_in_payload_111_imag;
      data_in_112_real <= io_data_in_payload_112_real;
      data_in_112_imag <= io_data_in_payload_112_imag;
      data_in_113_real <= io_data_in_payload_113_real;
      data_in_113_imag <= io_data_in_payload_113_imag;
      data_in_114_real <= io_data_in_payload_114_real;
      data_in_114_imag <= io_data_in_payload_114_imag;
      data_in_115_real <= io_data_in_payload_115_real;
      data_in_115_imag <= io_data_in_payload_115_imag;
      data_in_116_real <= io_data_in_payload_116_real;
      data_in_116_imag <= io_data_in_payload_116_imag;
      data_in_117_real <= io_data_in_payload_117_real;
      data_in_117_imag <= io_data_in_payload_117_imag;
      data_in_118_real <= io_data_in_payload_118_real;
      data_in_118_imag <= io_data_in_payload_118_imag;
      data_in_119_real <= io_data_in_payload_119_real;
      data_in_119_imag <= io_data_in_payload_119_imag;
      data_in_120_real <= io_data_in_payload_120_real;
      data_in_120_imag <= io_data_in_payload_120_imag;
      data_in_121_real <= io_data_in_payload_121_real;
      data_in_121_imag <= io_data_in_payload_121_imag;
      data_in_122_real <= io_data_in_payload_122_real;
      data_in_122_imag <= io_data_in_payload_122_imag;
      data_in_123_real <= io_data_in_payload_123_real;
      data_in_123_imag <= io_data_in_payload_123_imag;
      data_in_124_real <= io_data_in_payload_124_real;
      data_in_124_imag <= io_data_in_payload_124_imag;
      data_in_125_real <= io_data_in_payload_125_real;
      data_in_125_imag <= io_data_in_payload_125_imag;
      data_in_126_real <= io_data_in_payload_126_real;
      data_in_126_imag <= io_data_in_payload_126_imag;
      data_in_127_real <= io_data_in_payload_127_real;
      data_in_127_imag <= io_data_in_payload_127_imag;
    end
    io_data_in_valid_regNext <= io_data_in_valid;
    if((current_level_cnt_value == 3'b000))begin
      data_mid_0_real <= data_reorder_0_real;
      data_mid_0_imag <= data_reorder_0_imag;
      data_mid_1_real <= data_reorder_1_real;
      data_mid_1_imag <= data_reorder_1_imag;
      data_mid_2_real <= data_reorder_2_real;
      data_mid_2_imag <= data_reorder_2_imag;
      data_mid_3_real <= data_reorder_3_real;
      data_mid_3_imag <= data_reorder_3_imag;
      data_mid_4_real <= data_reorder_4_real;
      data_mid_4_imag <= data_reorder_4_imag;
      data_mid_5_real <= data_reorder_5_real;
      data_mid_5_imag <= data_reorder_5_imag;
      data_mid_6_real <= data_reorder_6_real;
      data_mid_6_imag <= data_reorder_6_imag;
      data_mid_7_real <= data_reorder_7_real;
      data_mid_7_imag <= data_reorder_7_imag;
      data_mid_8_real <= data_reorder_8_real;
      data_mid_8_imag <= data_reorder_8_imag;
      data_mid_9_real <= data_reorder_9_real;
      data_mid_9_imag <= data_reorder_9_imag;
      data_mid_10_real <= data_reorder_10_real;
      data_mid_10_imag <= data_reorder_10_imag;
      data_mid_11_real <= data_reorder_11_real;
      data_mid_11_imag <= data_reorder_11_imag;
      data_mid_12_real <= data_reorder_12_real;
      data_mid_12_imag <= data_reorder_12_imag;
      data_mid_13_real <= data_reorder_13_real;
      data_mid_13_imag <= data_reorder_13_imag;
      data_mid_14_real <= data_reorder_14_real;
      data_mid_14_imag <= data_reorder_14_imag;
      data_mid_15_real <= data_reorder_15_real;
      data_mid_15_imag <= data_reorder_15_imag;
      data_mid_16_real <= data_reorder_16_real;
      data_mid_16_imag <= data_reorder_16_imag;
      data_mid_17_real <= data_reorder_17_real;
      data_mid_17_imag <= data_reorder_17_imag;
      data_mid_18_real <= data_reorder_18_real;
      data_mid_18_imag <= data_reorder_18_imag;
      data_mid_19_real <= data_reorder_19_real;
      data_mid_19_imag <= data_reorder_19_imag;
      data_mid_20_real <= data_reorder_20_real;
      data_mid_20_imag <= data_reorder_20_imag;
      data_mid_21_real <= data_reorder_21_real;
      data_mid_21_imag <= data_reorder_21_imag;
      data_mid_22_real <= data_reorder_22_real;
      data_mid_22_imag <= data_reorder_22_imag;
      data_mid_23_real <= data_reorder_23_real;
      data_mid_23_imag <= data_reorder_23_imag;
      data_mid_24_real <= data_reorder_24_real;
      data_mid_24_imag <= data_reorder_24_imag;
      data_mid_25_real <= data_reorder_25_real;
      data_mid_25_imag <= data_reorder_25_imag;
      data_mid_26_real <= data_reorder_26_real;
      data_mid_26_imag <= data_reorder_26_imag;
      data_mid_27_real <= data_reorder_27_real;
      data_mid_27_imag <= data_reorder_27_imag;
      data_mid_28_real <= data_reorder_28_real;
      data_mid_28_imag <= data_reorder_28_imag;
      data_mid_29_real <= data_reorder_29_real;
      data_mid_29_imag <= data_reorder_29_imag;
      data_mid_30_real <= data_reorder_30_real;
      data_mid_30_imag <= data_reorder_30_imag;
      data_mid_31_real <= data_reorder_31_real;
      data_mid_31_imag <= data_reorder_31_imag;
      data_mid_32_real <= data_reorder_32_real;
      data_mid_32_imag <= data_reorder_32_imag;
      data_mid_33_real <= data_reorder_33_real;
      data_mid_33_imag <= data_reorder_33_imag;
      data_mid_34_real <= data_reorder_34_real;
      data_mid_34_imag <= data_reorder_34_imag;
      data_mid_35_real <= data_reorder_35_real;
      data_mid_35_imag <= data_reorder_35_imag;
      data_mid_36_real <= data_reorder_36_real;
      data_mid_36_imag <= data_reorder_36_imag;
      data_mid_37_real <= data_reorder_37_real;
      data_mid_37_imag <= data_reorder_37_imag;
      data_mid_38_real <= data_reorder_38_real;
      data_mid_38_imag <= data_reorder_38_imag;
      data_mid_39_real <= data_reorder_39_real;
      data_mid_39_imag <= data_reorder_39_imag;
      data_mid_40_real <= data_reorder_40_real;
      data_mid_40_imag <= data_reorder_40_imag;
      data_mid_41_real <= data_reorder_41_real;
      data_mid_41_imag <= data_reorder_41_imag;
      data_mid_42_real <= data_reorder_42_real;
      data_mid_42_imag <= data_reorder_42_imag;
      data_mid_43_real <= data_reorder_43_real;
      data_mid_43_imag <= data_reorder_43_imag;
      data_mid_44_real <= data_reorder_44_real;
      data_mid_44_imag <= data_reorder_44_imag;
      data_mid_45_real <= data_reorder_45_real;
      data_mid_45_imag <= data_reorder_45_imag;
      data_mid_46_real <= data_reorder_46_real;
      data_mid_46_imag <= data_reorder_46_imag;
      data_mid_47_real <= data_reorder_47_real;
      data_mid_47_imag <= data_reorder_47_imag;
      data_mid_48_real <= data_reorder_48_real;
      data_mid_48_imag <= data_reorder_48_imag;
      data_mid_49_real <= data_reorder_49_real;
      data_mid_49_imag <= data_reorder_49_imag;
      data_mid_50_real <= data_reorder_50_real;
      data_mid_50_imag <= data_reorder_50_imag;
      data_mid_51_real <= data_reorder_51_real;
      data_mid_51_imag <= data_reorder_51_imag;
      data_mid_52_real <= data_reorder_52_real;
      data_mid_52_imag <= data_reorder_52_imag;
      data_mid_53_real <= data_reorder_53_real;
      data_mid_53_imag <= data_reorder_53_imag;
      data_mid_54_real <= data_reorder_54_real;
      data_mid_54_imag <= data_reorder_54_imag;
      data_mid_55_real <= data_reorder_55_real;
      data_mid_55_imag <= data_reorder_55_imag;
      data_mid_56_real <= data_reorder_56_real;
      data_mid_56_imag <= data_reorder_56_imag;
      data_mid_57_real <= data_reorder_57_real;
      data_mid_57_imag <= data_reorder_57_imag;
      data_mid_58_real <= data_reorder_58_real;
      data_mid_58_imag <= data_reorder_58_imag;
      data_mid_59_real <= data_reorder_59_real;
      data_mid_59_imag <= data_reorder_59_imag;
      data_mid_60_real <= data_reorder_60_real;
      data_mid_60_imag <= data_reorder_60_imag;
      data_mid_61_real <= data_reorder_61_real;
      data_mid_61_imag <= data_reorder_61_imag;
      data_mid_62_real <= data_reorder_62_real;
      data_mid_62_imag <= data_reorder_62_imag;
      data_mid_63_real <= data_reorder_63_real;
      data_mid_63_imag <= data_reorder_63_imag;
      data_mid_64_real <= data_reorder_64_real;
      data_mid_64_imag <= data_reorder_64_imag;
      data_mid_65_real <= data_reorder_65_real;
      data_mid_65_imag <= data_reorder_65_imag;
      data_mid_66_real <= data_reorder_66_real;
      data_mid_66_imag <= data_reorder_66_imag;
      data_mid_67_real <= data_reorder_67_real;
      data_mid_67_imag <= data_reorder_67_imag;
      data_mid_68_real <= data_reorder_68_real;
      data_mid_68_imag <= data_reorder_68_imag;
      data_mid_69_real <= data_reorder_69_real;
      data_mid_69_imag <= data_reorder_69_imag;
      data_mid_70_real <= data_reorder_70_real;
      data_mid_70_imag <= data_reorder_70_imag;
      data_mid_71_real <= data_reorder_71_real;
      data_mid_71_imag <= data_reorder_71_imag;
      data_mid_72_real <= data_reorder_72_real;
      data_mid_72_imag <= data_reorder_72_imag;
      data_mid_73_real <= data_reorder_73_real;
      data_mid_73_imag <= data_reorder_73_imag;
      data_mid_74_real <= data_reorder_74_real;
      data_mid_74_imag <= data_reorder_74_imag;
      data_mid_75_real <= data_reorder_75_real;
      data_mid_75_imag <= data_reorder_75_imag;
      data_mid_76_real <= data_reorder_76_real;
      data_mid_76_imag <= data_reorder_76_imag;
      data_mid_77_real <= data_reorder_77_real;
      data_mid_77_imag <= data_reorder_77_imag;
      data_mid_78_real <= data_reorder_78_real;
      data_mid_78_imag <= data_reorder_78_imag;
      data_mid_79_real <= data_reorder_79_real;
      data_mid_79_imag <= data_reorder_79_imag;
      data_mid_80_real <= data_reorder_80_real;
      data_mid_80_imag <= data_reorder_80_imag;
      data_mid_81_real <= data_reorder_81_real;
      data_mid_81_imag <= data_reorder_81_imag;
      data_mid_82_real <= data_reorder_82_real;
      data_mid_82_imag <= data_reorder_82_imag;
      data_mid_83_real <= data_reorder_83_real;
      data_mid_83_imag <= data_reorder_83_imag;
      data_mid_84_real <= data_reorder_84_real;
      data_mid_84_imag <= data_reorder_84_imag;
      data_mid_85_real <= data_reorder_85_real;
      data_mid_85_imag <= data_reorder_85_imag;
      data_mid_86_real <= data_reorder_86_real;
      data_mid_86_imag <= data_reorder_86_imag;
      data_mid_87_real <= data_reorder_87_real;
      data_mid_87_imag <= data_reorder_87_imag;
      data_mid_88_real <= data_reorder_88_real;
      data_mid_88_imag <= data_reorder_88_imag;
      data_mid_89_real <= data_reorder_89_real;
      data_mid_89_imag <= data_reorder_89_imag;
      data_mid_90_real <= data_reorder_90_real;
      data_mid_90_imag <= data_reorder_90_imag;
      data_mid_91_real <= data_reorder_91_real;
      data_mid_91_imag <= data_reorder_91_imag;
      data_mid_92_real <= data_reorder_92_real;
      data_mid_92_imag <= data_reorder_92_imag;
      data_mid_93_real <= data_reorder_93_real;
      data_mid_93_imag <= data_reorder_93_imag;
      data_mid_94_real <= data_reorder_94_real;
      data_mid_94_imag <= data_reorder_94_imag;
      data_mid_95_real <= data_reorder_95_real;
      data_mid_95_imag <= data_reorder_95_imag;
      data_mid_96_real <= data_reorder_96_real;
      data_mid_96_imag <= data_reorder_96_imag;
      data_mid_97_real <= data_reorder_97_real;
      data_mid_97_imag <= data_reorder_97_imag;
      data_mid_98_real <= data_reorder_98_real;
      data_mid_98_imag <= data_reorder_98_imag;
      data_mid_99_real <= data_reorder_99_real;
      data_mid_99_imag <= data_reorder_99_imag;
      data_mid_100_real <= data_reorder_100_real;
      data_mid_100_imag <= data_reorder_100_imag;
      data_mid_101_real <= data_reorder_101_real;
      data_mid_101_imag <= data_reorder_101_imag;
      data_mid_102_real <= data_reorder_102_real;
      data_mid_102_imag <= data_reorder_102_imag;
      data_mid_103_real <= data_reorder_103_real;
      data_mid_103_imag <= data_reorder_103_imag;
      data_mid_104_real <= data_reorder_104_real;
      data_mid_104_imag <= data_reorder_104_imag;
      data_mid_105_real <= data_reorder_105_real;
      data_mid_105_imag <= data_reorder_105_imag;
      data_mid_106_real <= data_reorder_106_real;
      data_mid_106_imag <= data_reorder_106_imag;
      data_mid_107_real <= data_reorder_107_real;
      data_mid_107_imag <= data_reorder_107_imag;
      data_mid_108_real <= data_reorder_108_real;
      data_mid_108_imag <= data_reorder_108_imag;
      data_mid_109_real <= data_reorder_109_real;
      data_mid_109_imag <= data_reorder_109_imag;
      data_mid_110_real <= data_reorder_110_real;
      data_mid_110_imag <= data_reorder_110_imag;
      data_mid_111_real <= data_reorder_111_real;
      data_mid_111_imag <= data_reorder_111_imag;
      data_mid_112_real <= data_reorder_112_real;
      data_mid_112_imag <= data_reorder_112_imag;
      data_mid_113_real <= data_reorder_113_real;
      data_mid_113_imag <= data_reorder_113_imag;
      data_mid_114_real <= data_reorder_114_real;
      data_mid_114_imag <= data_reorder_114_imag;
      data_mid_115_real <= data_reorder_115_real;
      data_mid_115_imag <= data_reorder_115_imag;
      data_mid_116_real <= data_reorder_116_real;
      data_mid_116_imag <= data_reorder_116_imag;
      data_mid_117_real <= data_reorder_117_real;
      data_mid_117_imag <= data_reorder_117_imag;
      data_mid_118_real <= data_reorder_118_real;
      data_mid_118_imag <= data_reorder_118_imag;
      data_mid_119_real <= data_reorder_119_real;
      data_mid_119_imag <= data_reorder_119_imag;
      data_mid_120_real <= data_reorder_120_real;
      data_mid_120_imag <= data_reorder_120_imag;
      data_mid_121_real <= data_reorder_121_real;
      data_mid_121_imag <= data_reorder_121_imag;
      data_mid_122_real <= data_reorder_122_real;
      data_mid_122_imag <= data_reorder_122_imag;
      data_mid_123_real <= data_reorder_123_real;
      data_mid_123_imag <= data_reorder_123_imag;
      data_mid_124_real <= data_reorder_124_real;
      data_mid_124_imag <= data_reorder_124_imag;
      data_mid_125_real <= data_reorder_125_real;
      data_mid_125_imag <= data_reorder_125_imag;
      data_mid_126_real <= data_reorder_126_real;
      data_mid_126_imag <= data_reorder_126_imag;
      data_mid_127_real <= data_reorder_127_real;
      data_mid_127_imag <= data_reorder_127_imag;
    end else begin
      if((current_level_cnt_value == 3'b001))begin
        data_mid_1_real <= _zz_2697[15 : 0];
        data_mid_1_imag <= _zz_2701[15 : 0];
        data_mid_0_real <= _zz_2705[15 : 0];
        data_mid_0_imag <= _zz_2709[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_3_real <= _zz_2719[15 : 0];
        data_mid_3_imag <= _zz_2723[15 : 0];
        data_mid_2_real <= _zz_2727[15 : 0];
        data_mid_2_imag <= _zz_2731[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_5_real <= _zz_2741[15 : 0];
        data_mid_5_imag <= _zz_2745[15 : 0];
        data_mid_4_real <= _zz_2749[15 : 0];
        data_mid_4_imag <= _zz_2753[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_7_real <= _zz_2763[15 : 0];
        data_mid_7_imag <= _zz_2767[15 : 0];
        data_mid_6_real <= _zz_2771[15 : 0];
        data_mid_6_imag <= _zz_2775[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_9_real <= _zz_2785[15 : 0];
        data_mid_9_imag <= _zz_2789[15 : 0];
        data_mid_8_real <= _zz_2793[15 : 0];
        data_mid_8_imag <= _zz_2797[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_11_real <= _zz_2807[15 : 0];
        data_mid_11_imag <= _zz_2811[15 : 0];
        data_mid_10_real <= _zz_2815[15 : 0];
        data_mid_10_imag <= _zz_2819[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_13_real <= _zz_2829[15 : 0];
        data_mid_13_imag <= _zz_2833[15 : 0];
        data_mid_12_real <= _zz_2837[15 : 0];
        data_mid_12_imag <= _zz_2841[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_15_real <= _zz_2851[15 : 0];
        data_mid_15_imag <= _zz_2855[15 : 0];
        data_mid_14_real <= _zz_2859[15 : 0];
        data_mid_14_imag <= _zz_2863[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_17_real <= _zz_2873[15 : 0];
        data_mid_17_imag <= _zz_2877[15 : 0];
        data_mid_16_real <= _zz_2881[15 : 0];
        data_mid_16_imag <= _zz_2885[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_19_real <= _zz_2895[15 : 0];
        data_mid_19_imag <= _zz_2899[15 : 0];
        data_mid_18_real <= _zz_2903[15 : 0];
        data_mid_18_imag <= _zz_2907[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_21_real <= _zz_2917[15 : 0];
        data_mid_21_imag <= _zz_2921[15 : 0];
        data_mid_20_real <= _zz_2925[15 : 0];
        data_mid_20_imag <= _zz_2929[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_23_real <= _zz_2939[15 : 0];
        data_mid_23_imag <= _zz_2943[15 : 0];
        data_mid_22_real <= _zz_2947[15 : 0];
        data_mid_22_imag <= _zz_2951[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_25_real <= _zz_2961[15 : 0];
        data_mid_25_imag <= _zz_2965[15 : 0];
        data_mid_24_real <= _zz_2969[15 : 0];
        data_mid_24_imag <= _zz_2973[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_27_real <= _zz_2983[15 : 0];
        data_mid_27_imag <= _zz_2987[15 : 0];
        data_mid_26_real <= _zz_2991[15 : 0];
        data_mid_26_imag <= _zz_2995[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_29_real <= _zz_3005[15 : 0];
        data_mid_29_imag <= _zz_3009[15 : 0];
        data_mid_28_real <= _zz_3013[15 : 0];
        data_mid_28_imag <= _zz_3017[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_31_real <= _zz_3027[15 : 0];
        data_mid_31_imag <= _zz_3031[15 : 0];
        data_mid_30_real <= _zz_3035[15 : 0];
        data_mid_30_imag <= _zz_3039[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_33_real <= _zz_3049[15 : 0];
        data_mid_33_imag <= _zz_3053[15 : 0];
        data_mid_32_real <= _zz_3057[15 : 0];
        data_mid_32_imag <= _zz_3061[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_35_real <= _zz_3071[15 : 0];
        data_mid_35_imag <= _zz_3075[15 : 0];
        data_mid_34_real <= _zz_3079[15 : 0];
        data_mid_34_imag <= _zz_3083[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_37_real <= _zz_3093[15 : 0];
        data_mid_37_imag <= _zz_3097[15 : 0];
        data_mid_36_real <= _zz_3101[15 : 0];
        data_mid_36_imag <= _zz_3105[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_39_real <= _zz_3115[15 : 0];
        data_mid_39_imag <= _zz_3119[15 : 0];
        data_mid_38_real <= _zz_3123[15 : 0];
        data_mid_38_imag <= _zz_3127[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_41_real <= _zz_3137[15 : 0];
        data_mid_41_imag <= _zz_3141[15 : 0];
        data_mid_40_real <= _zz_3145[15 : 0];
        data_mid_40_imag <= _zz_3149[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_43_real <= _zz_3159[15 : 0];
        data_mid_43_imag <= _zz_3163[15 : 0];
        data_mid_42_real <= _zz_3167[15 : 0];
        data_mid_42_imag <= _zz_3171[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_45_real <= _zz_3181[15 : 0];
        data_mid_45_imag <= _zz_3185[15 : 0];
        data_mid_44_real <= _zz_3189[15 : 0];
        data_mid_44_imag <= _zz_3193[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_47_real <= _zz_3203[15 : 0];
        data_mid_47_imag <= _zz_3207[15 : 0];
        data_mid_46_real <= _zz_3211[15 : 0];
        data_mid_46_imag <= _zz_3215[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_49_real <= _zz_3225[15 : 0];
        data_mid_49_imag <= _zz_3229[15 : 0];
        data_mid_48_real <= _zz_3233[15 : 0];
        data_mid_48_imag <= _zz_3237[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_51_real <= _zz_3247[15 : 0];
        data_mid_51_imag <= _zz_3251[15 : 0];
        data_mid_50_real <= _zz_3255[15 : 0];
        data_mid_50_imag <= _zz_3259[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_53_real <= _zz_3269[15 : 0];
        data_mid_53_imag <= _zz_3273[15 : 0];
        data_mid_52_real <= _zz_3277[15 : 0];
        data_mid_52_imag <= _zz_3281[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_55_real <= _zz_3291[15 : 0];
        data_mid_55_imag <= _zz_3295[15 : 0];
        data_mid_54_real <= _zz_3299[15 : 0];
        data_mid_54_imag <= _zz_3303[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_57_real <= _zz_3313[15 : 0];
        data_mid_57_imag <= _zz_3317[15 : 0];
        data_mid_56_real <= _zz_3321[15 : 0];
        data_mid_56_imag <= _zz_3325[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_59_real <= _zz_3335[15 : 0];
        data_mid_59_imag <= _zz_3339[15 : 0];
        data_mid_58_real <= _zz_3343[15 : 0];
        data_mid_58_imag <= _zz_3347[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_61_real <= _zz_3357[15 : 0];
        data_mid_61_imag <= _zz_3361[15 : 0];
        data_mid_60_real <= _zz_3365[15 : 0];
        data_mid_60_imag <= _zz_3369[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_63_real <= _zz_3379[15 : 0];
        data_mid_63_imag <= _zz_3383[15 : 0];
        data_mid_62_real <= _zz_3387[15 : 0];
        data_mid_62_imag <= _zz_3391[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_65_real <= _zz_3401[15 : 0];
        data_mid_65_imag <= _zz_3405[15 : 0];
        data_mid_64_real <= _zz_3409[15 : 0];
        data_mid_64_imag <= _zz_3413[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_67_real <= _zz_3423[15 : 0];
        data_mid_67_imag <= _zz_3427[15 : 0];
        data_mid_66_real <= _zz_3431[15 : 0];
        data_mid_66_imag <= _zz_3435[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_69_real <= _zz_3445[15 : 0];
        data_mid_69_imag <= _zz_3449[15 : 0];
        data_mid_68_real <= _zz_3453[15 : 0];
        data_mid_68_imag <= _zz_3457[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_71_real <= _zz_3467[15 : 0];
        data_mid_71_imag <= _zz_3471[15 : 0];
        data_mid_70_real <= _zz_3475[15 : 0];
        data_mid_70_imag <= _zz_3479[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_73_real <= _zz_3489[15 : 0];
        data_mid_73_imag <= _zz_3493[15 : 0];
        data_mid_72_real <= _zz_3497[15 : 0];
        data_mid_72_imag <= _zz_3501[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_75_real <= _zz_3511[15 : 0];
        data_mid_75_imag <= _zz_3515[15 : 0];
        data_mid_74_real <= _zz_3519[15 : 0];
        data_mid_74_imag <= _zz_3523[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_77_real <= _zz_3533[15 : 0];
        data_mid_77_imag <= _zz_3537[15 : 0];
        data_mid_76_real <= _zz_3541[15 : 0];
        data_mid_76_imag <= _zz_3545[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_79_real <= _zz_3555[15 : 0];
        data_mid_79_imag <= _zz_3559[15 : 0];
        data_mid_78_real <= _zz_3563[15 : 0];
        data_mid_78_imag <= _zz_3567[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_81_real <= _zz_3577[15 : 0];
        data_mid_81_imag <= _zz_3581[15 : 0];
        data_mid_80_real <= _zz_3585[15 : 0];
        data_mid_80_imag <= _zz_3589[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_83_real <= _zz_3599[15 : 0];
        data_mid_83_imag <= _zz_3603[15 : 0];
        data_mid_82_real <= _zz_3607[15 : 0];
        data_mid_82_imag <= _zz_3611[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_85_real <= _zz_3621[15 : 0];
        data_mid_85_imag <= _zz_3625[15 : 0];
        data_mid_84_real <= _zz_3629[15 : 0];
        data_mid_84_imag <= _zz_3633[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_87_real <= _zz_3643[15 : 0];
        data_mid_87_imag <= _zz_3647[15 : 0];
        data_mid_86_real <= _zz_3651[15 : 0];
        data_mid_86_imag <= _zz_3655[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_89_real <= _zz_3665[15 : 0];
        data_mid_89_imag <= _zz_3669[15 : 0];
        data_mid_88_real <= _zz_3673[15 : 0];
        data_mid_88_imag <= _zz_3677[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_91_real <= _zz_3687[15 : 0];
        data_mid_91_imag <= _zz_3691[15 : 0];
        data_mid_90_real <= _zz_3695[15 : 0];
        data_mid_90_imag <= _zz_3699[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_93_real <= _zz_3709[15 : 0];
        data_mid_93_imag <= _zz_3713[15 : 0];
        data_mid_92_real <= _zz_3717[15 : 0];
        data_mid_92_imag <= _zz_3721[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_95_real <= _zz_3731[15 : 0];
        data_mid_95_imag <= _zz_3735[15 : 0];
        data_mid_94_real <= _zz_3739[15 : 0];
        data_mid_94_imag <= _zz_3743[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_97_real <= _zz_3753[15 : 0];
        data_mid_97_imag <= _zz_3757[15 : 0];
        data_mid_96_real <= _zz_3761[15 : 0];
        data_mid_96_imag <= _zz_3765[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_99_real <= _zz_3775[15 : 0];
        data_mid_99_imag <= _zz_3779[15 : 0];
        data_mid_98_real <= _zz_3783[15 : 0];
        data_mid_98_imag <= _zz_3787[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_101_real <= _zz_3797[15 : 0];
        data_mid_101_imag <= _zz_3801[15 : 0];
        data_mid_100_real <= _zz_3805[15 : 0];
        data_mid_100_imag <= _zz_3809[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_103_real <= _zz_3819[15 : 0];
        data_mid_103_imag <= _zz_3823[15 : 0];
        data_mid_102_real <= _zz_3827[15 : 0];
        data_mid_102_imag <= _zz_3831[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_105_real <= _zz_3841[15 : 0];
        data_mid_105_imag <= _zz_3845[15 : 0];
        data_mid_104_real <= _zz_3849[15 : 0];
        data_mid_104_imag <= _zz_3853[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_107_real <= _zz_3863[15 : 0];
        data_mid_107_imag <= _zz_3867[15 : 0];
        data_mid_106_real <= _zz_3871[15 : 0];
        data_mid_106_imag <= _zz_3875[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_109_real <= _zz_3885[15 : 0];
        data_mid_109_imag <= _zz_3889[15 : 0];
        data_mid_108_real <= _zz_3893[15 : 0];
        data_mid_108_imag <= _zz_3897[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_111_real <= _zz_3907[15 : 0];
        data_mid_111_imag <= _zz_3911[15 : 0];
        data_mid_110_real <= _zz_3915[15 : 0];
        data_mid_110_imag <= _zz_3919[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_113_real <= _zz_3929[15 : 0];
        data_mid_113_imag <= _zz_3933[15 : 0];
        data_mid_112_real <= _zz_3937[15 : 0];
        data_mid_112_imag <= _zz_3941[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_115_real <= _zz_3951[15 : 0];
        data_mid_115_imag <= _zz_3955[15 : 0];
        data_mid_114_real <= _zz_3959[15 : 0];
        data_mid_114_imag <= _zz_3963[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_117_real <= _zz_3973[15 : 0];
        data_mid_117_imag <= _zz_3977[15 : 0];
        data_mid_116_real <= _zz_3981[15 : 0];
        data_mid_116_imag <= _zz_3985[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_119_real <= _zz_3995[15 : 0];
        data_mid_119_imag <= _zz_3999[15 : 0];
        data_mid_118_real <= _zz_4003[15 : 0];
        data_mid_118_imag <= _zz_4007[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_121_real <= _zz_4017[15 : 0];
        data_mid_121_imag <= _zz_4021[15 : 0];
        data_mid_120_real <= _zz_4025[15 : 0];
        data_mid_120_imag <= _zz_4029[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_123_real <= _zz_4039[15 : 0];
        data_mid_123_imag <= _zz_4043[15 : 0];
        data_mid_122_real <= _zz_4047[15 : 0];
        data_mid_122_imag <= _zz_4051[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_125_real <= _zz_4061[15 : 0];
        data_mid_125_imag <= _zz_4065[15 : 0];
        data_mid_124_real <= _zz_4069[15 : 0];
        data_mid_124_imag <= _zz_4073[15 : 0];
      end
      if((current_level_cnt_value == 3'b001))begin
        data_mid_127_real <= _zz_4083[15 : 0];
        data_mid_127_imag <= _zz_4087[15 : 0];
        data_mid_126_real <= _zz_4091[15 : 0];
        data_mid_126_imag <= _zz_4095[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_2_real <= _zz_4105[15 : 0];
        data_mid_2_imag <= _zz_4109[15 : 0];
        data_mid_0_real <= _zz_4113[15 : 0];
        data_mid_0_imag <= _zz_4117[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_3_real <= _zz_4127[15 : 0];
        data_mid_3_imag <= _zz_4131[15 : 0];
        data_mid_1_real <= _zz_4135[15 : 0];
        data_mid_1_imag <= _zz_4139[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_6_real <= _zz_4149[15 : 0];
        data_mid_6_imag <= _zz_4153[15 : 0];
        data_mid_4_real <= _zz_4157[15 : 0];
        data_mid_4_imag <= _zz_4161[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_7_real <= _zz_4171[15 : 0];
        data_mid_7_imag <= _zz_4175[15 : 0];
        data_mid_5_real <= _zz_4179[15 : 0];
        data_mid_5_imag <= _zz_4183[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_10_real <= _zz_4193[15 : 0];
        data_mid_10_imag <= _zz_4197[15 : 0];
        data_mid_8_real <= _zz_4201[15 : 0];
        data_mid_8_imag <= _zz_4205[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_11_real <= _zz_4215[15 : 0];
        data_mid_11_imag <= _zz_4219[15 : 0];
        data_mid_9_real <= _zz_4223[15 : 0];
        data_mid_9_imag <= _zz_4227[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_14_real <= _zz_4237[15 : 0];
        data_mid_14_imag <= _zz_4241[15 : 0];
        data_mid_12_real <= _zz_4245[15 : 0];
        data_mid_12_imag <= _zz_4249[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_15_real <= _zz_4259[15 : 0];
        data_mid_15_imag <= _zz_4263[15 : 0];
        data_mid_13_real <= _zz_4267[15 : 0];
        data_mid_13_imag <= _zz_4271[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_18_real <= _zz_4281[15 : 0];
        data_mid_18_imag <= _zz_4285[15 : 0];
        data_mid_16_real <= _zz_4289[15 : 0];
        data_mid_16_imag <= _zz_4293[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_19_real <= _zz_4303[15 : 0];
        data_mid_19_imag <= _zz_4307[15 : 0];
        data_mid_17_real <= _zz_4311[15 : 0];
        data_mid_17_imag <= _zz_4315[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_22_real <= _zz_4325[15 : 0];
        data_mid_22_imag <= _zz_4329[15 : 0];
        data_mid_20_real <= _zz_4333[15 : 0];
        data_mid_20_imag <= _zz_4337[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_23_real <= _zz_4347[15 : 0];
        data_mid_23_imag <= _zz_4351[15 : 0];
        data_mid_21_real <= _zz_4355[15 : 0];
        data_mid_21_imag <= _zz_4359[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_26_real <= _zz_4369[15 : 0];
        data_mid_26_imag <= _zz_4373[15 : 0];
        data_mid_24_real <= _zz_4377[15 : 0];
        data_mid_24_imag <= _zz_4381[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_27_real <= _zz_4391[15 : 0];
        data_mid_27_imag <= _zz_4395[15 : 0];
        data_mid_25_real <= _zz_4399[15 : 0];
        data_mid_25_imag <= _zz_4403[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_30_real <= _zz_4413[15 : 0];
        data_mid_30_imag <= _zz_4417[15 : 0];
        data_mid_28_real <= _zz_4421[15 : 0];
        data_mid_28_imag <= _zz_4425[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_31_real <= _zz_4435[15 : 0];
        data_mid_31_imag <= _zz_4439[15 : 0];
        data_mid_29_real <= _zz_4443[15 : 0];
        data_mid_29_imag <= _zz_4447[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_34_real <= _zz_4457[15 : 0];
        data_mid_34_imag <= _zz_4461[15 : 0];
        data_mid_32_real <= _zz_4465[15 : 0];
        data_mid_32_imag <= _zz_4469[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_35_real <= _zz_4479[15 : 0];
        data_mid_35_imag <= _zz_4483[15 : 0];
        data_mid_33_real <= _zz_4487[15 : 0];
        data_mid_33_imag <= _zz_4491[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_38_real <= _zz_4501[15 : 0];
        data_mid_38_imag <= _zz_4505[15 : 0];
        data_mid_36_real <= _zz_4509[15 : 0];
        data_mid_36_imag <= _zz_4513[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_39_real <= _zz_4523[15 : 0];
        data_mid_39_imag <= _zz_4527[15 : 0];
        data_mid_37_real <= _zz_4531[15 : 0];
        data_mid_37_imag <= _zz_4535[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_42_real <= _zz_4545[15 : 0];
        data_mid_42_imag <= _zz_4549[15 : 0];
        data_mid_40_real <= _zz_4553[15 : 0];
        data_mid_40_imag <= _zz_4557[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_43_real <= _zz_4567[15 : 0];
        data_mid_43_imag <= _zz_4571[15 : 0];
        data_mid_41_real <= _zz_4575[15 : 0];
        data_mid_41_imag <= _zz_4579[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_46_real <= _zz_4589[15 : 0];
        data_mid_46_imag <= _zz_4593[15 : 0];
        data_mid_44_real <= _zz_4597[15 : 0];
        data_mid_44_imag <= _zz_4601[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_47_real <= _zz_4611[15 : 0];
        data_mid_47_imag <= _zz_4615[15 : 0];
        data_mid_45_real <= _zz_4619[15 : 0];
        data_mid_45_imag <= _zz_4623[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_50_real <= _zz_4633[15 : 0];
        data_mid_50_imag <= _zz_4637[15 : 0];
        data_mid_48_real <= _zz_4641[15 : 0];
        data_mid_48_imag <= _zz_4645[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_51_real <= _zz_4655[15 : 0];
        data_mid_51_imag <= _zz_4659[15 : 0];
        data_mid_49_real <= _zz_4663[15 : 0];
        data_mid_49_imag <= _zz_4667[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_54_real <= _zz_4677[15 : 0];
        data_mid_54_imag <= _zz_4681[15 : 0];
        data_mid_52_real <= _zz_4685[15 : 0];
        data_mid_52_imag <= _zz_4689[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_55_real <= _zz_4699[15 : 0];
        data_mid_55_imag <= _zz_4703[15 : 0];
        data_mid_53_real <= _zz_4707[15 : 0];
        data_mid_53_imag <= _zz_4711[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_58_real <= _zz_4721[15 : 0];
        data_mid_58_imag <= _zz_4725[15 : 0];
        data_mid_56_real <= _zz_4729[15 : 0];
        data_mid_56_imag <= _zz_4733[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_59_real <= _zz_4743[15 : 0];
        data_mid_59_imag <= _zz_4747[15 : 0];
        data_mid_57_real <= _zz_4751[15 : 0];
        data_mid_57_imag <= _zz_4755[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_62_real <= _zz_4765[15 : 0];
        data_mid_62_imag <= _zz_4769[15 : 0];
        data_mid_60_real <= _zz_4773[15 : 0];
        data_mid_60_imag <= _zz_4777[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_63_real <= _zz_4787[15 : 0];
        data_mid_63_imag <= _zz_4791[15 : 0];
        data_mid_61_real <= _zz_4795[15 : 0];
        data_mid_61_imag <= _zz_4799[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_66_real <= _zz_4809[15 : 0];
        data_mid_66_imag <= _zz_4813[15 : 0];
        data_mid_64_real <= _zz_4817[15 : 0];
        data_mid_64_imag <= _zz_4821[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_67_real <= _zz_4831[15 : 0];
        data_mid_67_imag <= _zz_4835[15 : 0];
        data_mid_65_real <= _zz_4839[15 : 0];
        data_mid_65_imag <= _zz_4843[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_70_real <= _zz_4853[15 : 0];
        data_mid_70_imag <= _zz_4857[15 : 0];
        data_mid_68_real <= _zz_4861[15 : 0];
        data_mid_68_imag <= _zz_4865[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_71_real <= _zz_4875[15 : 0];
        data_mid_71_imag <= _zz_4879[15 : 0];
        data_mid_69_real <= _zz_4883[15 : 0];
        data_mid_69_imag <= _zz_4887[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_74_real <= _zz_4897[15 : 0];
        data_mid_74_imag <= _zz_4901[15 : 0];
        data_mid_72_real <= _zz_4905[15 : 0];
        data_mid_72_imag <= _zz_4909[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_75_real <= _zz_4919[15 : 0];
        data_mid_75_imag <= _zz_4923[15 : 0];
        data_mid_73_real <= _zz_4927[15 : 0];
        data_mid_73_imag <= _zz_4931[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_78_real <= _zz_4941[15 : 0];
        data_mid_78_imag <= _zz_4945[15 : 0];
        data_mid_76_real <= _zz_4949[15 : 0];
        data_mid_76_imag <= _zz_4953[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_79_real <= _zz_4963[15 : 0];
        data_mid_79_imag <= _zz_4967[15 : 0];
        data_mid_77_real <= _zz_4971[15 : 0];
        data_mid_77_imag <= _zz_4975[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_82_real <= _zz_4985[15 : 0];
        data_mid_82_imag <= _zz_4989[15 : 0];
        data_mid_80_real <= _zz_4993[15 : 0];
        data_mid_80_imag <= _zz_4997[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_83_real <= _zz_5007[15 : 0];
        data_mid_83_imag <= _zz_5011[15 : 0];
        data_mid_81_real <= _zz_5015[15 : 0];
        data_mid_81_imag <= _zz_5019[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_86_real <= _zz_5029[15 : 0];
        data_mid_86_imag <= _zz_5033[15 : 0];
        data_mid_84_real <= _zz_5037[15 : 0];
        data_mid_84_imag <= _zz_5041[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_87_real <= _zz_5051[15 : 0];
        data_mid_87_imag <= _zz_5055[15 : 0];
        data_mid_85_real <= _zz_5059[15 : 0];
        data_mid_85_imag <= _zz_5063[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_90_real <= _zz_5073[15 : 0];
        data_mid_90_imag <= _zz_5077[15 : 0];
        data_mid_88_real <= _zz_5081[15 : 0];
        data_mid_88_imag <= _zz_5085[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_91_real <= _zz_5095[15 : 0];
        data_mid_91_imag <= _zz_5099[15 : 0];
        data_mid_89_real <= _zz_5103[15 : 0];
        data_mid_89_imag <= _zz_5107[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_94_real <= _zz_5117[15 : 0];
        data_mid_94_imag <= _zz_5121[15 : 0];
        data_mid_92_real <= _zz_5125[15 : 0];
        data_mid_92_imag <= _zz_5129[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_95_real <= _zz_5139[15 : 0];
        data_mid_95_imag <= _zz_5143[15 : 0];
        data_mid_93_real <= _zz_5147[15 : 0];
        data_mid_93_imag <= _zz_5151[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_98_real <= _zz_5161[15 : 0];
        data_mid_98_imag <= _zz_5165[15 : 0];
        data_mid_96_real <= _zz_5169[15 : 0];
        data_mid_96_imag <= _zz_5173[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_99_real <= _zz_5183[15 : 0];
        data_mid_99_imag <= _zz_5187[15 : 0];
        data_mid_97_real <= _zz_5191[15 : 0];
        data_mid_97_imag <= _zz_5195[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_102_real <= _zz_5205[15 : 0];
        data_mid_102_imag <= _zz_5209[15 : 0];
        data_mid_100_real <= _zz_5213[15 : 0];
        data_mid_100_imag <= _zz_5217[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_103_real <= _zz_5227[15 : 0];
        data_mid_103_imag <= _zz_5231[15 : 0];
        data_mid_101_real <= _zz_5235[15 : 0];
        data_mid_101_imag <= _zz_5239[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_106_real <= _zz_5249[15 : 0];
        data_mid_106_imag <= _zz_5253[15 : 0];
        data_mid_104_real <= _zz_5257[15 : 0];
        data_mid_104_imag <= _zz_5261[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_107_real <= _zz_5271[15 : 0];
        data_mid_107_imag <= _zz_5275[15 : 0];
        data_mid_105_real <= _zz_5279[15 : 0];
        data_mid_105_imag <= _zz_5283[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_110_real <= _zz_5293[15 : 0];
        data_mid_110_imag <= _zz_5297[15 : 0];
        data_mid_108_real <= _zz_5301[15 : 0];
        data_mid_108_imag <= _zz_5305[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_111_real <= _zz_5315[15 : 0];
        data_mid_111_imag <= _zz_5319[15 : 0];
        data_mid_109_real <= _zz_5323[15 : 0];
        data_mid_109_imag <= _zz_5327[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_114_real <= _zz_5337[15 : 0];
        data_mid_114_imag <= _zz_5341[15 : 0];
        data_mid_112_real <= _zz_5345[15 : 0];
        data_mid_112_imag <= _zz_5349[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_115_real <= _zz_5359[15 : 0];
        data_mid_115_imag <= _zz_5363[15 : 0];
        data_mid_113_real <= _zz_5367[15 : 0];
        data_mid_113_imag <= _zz_5371[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_118_real <= _zz_5381[15 : 0];
        data_mid_118_imag <= _zz_5385[15 : 0];
        data_mid_116_real <= _zz_5389[15 : 0];
        data_mid_116_imag <= _zz_5393[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_119_real <= _zz_5403[15 : 0];
        data_mid_119_imag <= _zz_5407[15 : 0];
        data_mid_117_real <= _zz_5411[15 : 0];
        data_mid_117_imag <= _zz_5415[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_122_real <= _zz_5425[15 : 0];
        data_mid_122_imag <= _zz_5429[15 : 0];
        data_mid_120_real <= _zz_5433[15 : 0];
        data_mid_120_imag <= _zz_5437[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_123_real <= _zz_5447[15 : 0];
        data_mid_123_imag <= _zz_5451[15 : 0];
        data_mid_121_real <= _zz_5455[15 : 0];
        data_mid_121_imag <= _zz_5459[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_126_real <= _zz_5469[15 : 0];
        data_mid_126_imag <= _zz_5473[15 : 0];
        data_mid_124_real <= _zz_5477[15 : 0];
        data_mid_124_imag <= _zz_5481[15 : 0];
      end
      if((current_level_cnt_value == 3'b010))begin
        data_mid_127_real <= _zz_5491[15 : 0];
        data_mid_127_imag <= _zz_5495[15 : 0];
        data_mid_125_real <= _zz_5499[15 : 0];
        data_mid_125_imag <= _zz_5503[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_4_real <= _zz_5513[15 : 0];
        data_mid_4_imag <= _zz_5517[15 : 0];
        data_mid_0_real <= _zz_5521[15 : 0];
        data_mid_0_imag <= _zz_5525[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_5_real <= _zz_5535[15 : 0];
        data_mid_5_imag <= _zz_5539[15 : 0];
        data_mid_1_real <= _zz_5543[15 : 0];
        data_mid_1_imag <= _zz_5547[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_6_real <= _zz_5557[15 : 0];
        data_mid_6_imag <= _zz_5561[15 : 0];
        data_mid_2_real <= _zz_5565[15 : 0];
        data_mid_2_imag <= _zz_5569[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_7_real <= _zz_5579[15 : 0];
        data_mid_7_imag <= _zz_5583[15 : 0];
        data_mid_3_real <= _zz_5587[15 : 0];
        data_mid_3_imag <= _zz_5591[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_12_real <= _zz_5601[15 : 0];
        data_mid_12_imag <= _zz_5605[15 : 0];
        data_mid_8_real <= _zz_5609[15 : 0];
        data_mid_8_imag <= _zz_5613[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_13_real <= _zz_5623[15 : 0];
        data_mid_13_imag <= _zz_5627[15 : 0];
        data_mid_9_real <= _zz_5631[15 : 0];
        data_mid_9_imag <= _zz_5635[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_14_real <= _zz_5645[15 : 0];
        data_mid_14_imag <= _zz_5649[15 : 0];
        data_mid_10_real <= _zz_5653[15 : 0];
        data_mid_10_imag <= _zz_5657[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_15_real <= _zz_5667[15 : 0];
        data_mid_15_imag <= _zz_5671[15 : 0];
        data_mid_11_real <= _zz_5675[15 : 0];
        data_mid_11_imag <= _zz_5679[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_20_real <= _zz_5689[15 : 0];
        data_mid_20_imag <= _zz_5693[15 : 0];
        data_mid_16_real <= _zz_5697[15 : 0];
        data_mid_16_imag <= _zz_5701[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_21_real <= _zz_5711[15 : 0];
        data_mid_21_imag <= _zz_5715[15 : 0];
        data_mid_17_real <= _zz_5719[15 : 0];
        data_mid_17_imag <= _zz_5723[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_22_real <= _zz_5733[15 : 0];
        data_mid_22_imag <= _zz_5737[15 : 0];
        data_mid_18_real <= _zz_5741[15 : 0];
        data_mid_18_imag <= _zz_5745[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_23_real <= _zz_5755[15 : 0];
        data_mid_23_imag <= _zz_5759[15 : 0];
        data_mid_19_real <= _zz_5763[15 : 0];
        data_mid_19_imag <= _zz_5767[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_28_real <= _zz_5777[15 : 0];
        data_mid_28_imag <= _zz_5781[15 : 0];
        data_mid_24_real <= _zz_5785[15 : 0];
        data_mid_24_imag <= _zz_5789[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_29_real <= _zz_5799[15 : 0];
        data_mid_29_imag <= _zz_5803[15 : 0];
        data_mid_25_real <= _zz_5807[15 : 0];
        data_mid_25_imag <= _zz_5811[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_30_real <= _zz_5821[15 : 0];
        data_mid_30_imag <= _zz_5825[15 : 0];
        data_mid_26_real <= _zz_5829[15 : 0];
        data_mid_26_imag <= _zz_5833[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_31_real <= _zz_5843[15 : 0];
        data_mid_31_imag <= _zz_5847[15 : 0];
        data_mid_27_real <= _zz_5851[15 : 0];
        data_mid_27_imag <= _zz_5855[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_36_real <= _zz_5865[15 : 0];
        data_mid_36_imag <= _zz_5869[15 : 0];
        data_mid_32_real <= _zz_5873[15 : 0];
        data_mid_32_imag <= _zz_5877[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_37_real <= _zz_5887[15 : 0];
        data_mid_37_imag <= _zz_5891[15 : 0];
        data_mid_33_real <= _zz_5895[15 : 0];
        data_mid_33_imag <= _zz_5899[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_38_real <= _zz_5909[15 : 0];
        data_mid_38_imag <= _zz_5913[15 : 0];
        data_mid_34_real <= _zz_5917[15 : 0];
        data_mid_34_imag <= _zz_5921[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_39_real <= _zz_5931[15 : 0];
        data_mid_39_imag <= _zz_5935[15 : 0];
        data_mid_35_real <= _zz_5939[15 : 0];
        data_mid_35_imag <= _zz_5943[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_44_real <= _zz_5953[15 : 0];
        data_mid_44_imag <= _zz_5957[15 : 0];
        data_mid_40_real <= _zz_5961[15 : 0];
        data_mid_40_imag <= _zz_5965[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_45_real <= _zz_5975[15 : 0];
        data_mid_45_imag <= _zz_5979[15 : 0];
        data_mid_41_real <= _zz_5983[15 : 0];
        data_mid_41_imag <= _zz_5987[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_46_real <= _zz_5997[15 : 0];
        data_mid_46_imag <= _zz_6001[15 : 0];
        data_mid_42_real <= _zz_6005[15 : 0];
        data_mid_42_imag <= _zz_6009[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_47_real <= _zz_6019[15 : 0];
        data_mid_47_imag <= _zz_6023[15 : 0];
        data_mid_43_real <= _zz_6027[15 : 0];
        data_mid_43_imag <= _zz_6031[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_52_real <= _zz_6041[15 : 0];
        data_mid_52_imag <= _zz_6045[15 : 0];
        data_mid_48_real <= _zz_6049[15 : 0];
        data_mid_48_imag <= _zz_6053[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_53_real <= _zz_6063[15 : 0];
        data_mid_53_imag <= _zz_6067[15 : 0];
        data_mid_49_real <= _zz_6071[15 : 0];
        data_mid_49_imag <= _zz_6075[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_54_real <= _zz_6085[15 : 0];
        data_mid_54_imag <= _zz_6089[15 : 0];
        data_mid_50_real <= _zz_6093[15 : 0];
        data_mid_50_imag <= _zz_6097[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_55_real <= _zz_6107[15 : 0];
        data_mid_55_imag <= _zz_6111[15 : 0];
        data_mid_51_real <= _zz_6115[15 : 0];
        data_mid_51_imag <= _zz_6119[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_60_real <= _zz_6129[15 : 0];
        data_mid_60_imag <= _zz_6133[15 : 0];
        data_mid_56_real <= _zz_6137[15 : 0];
        data_mid_56_imag <= _zz_6141[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_61_real <= _zz_6151[15 : 0];
        data_mid_61_imag <= _zz_6155[15 : 0];
        data_mid_57_real <= _zz_6159[15 : 0];
        data_mid_57_imag <= _zz_6163[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_62_real <= _zz_6173[15 : 0];
        data_mid_62_imag <= _zz_6177[15 : 0];
        data_mid_58_real <= _zz_6181[15 : 0];
        data_mid_58_imag <= _zz_6185[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_63_real <= _zz_6195[15 : 0];
        data_mid_63_imag <= _zz_6199[15 : 0];
        data_mid_59_real <= _zz_6203[15 : 0];
        data_mid_59_imag <= _zz_6207[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_68_real <= _zz_6217[15 : 0];
        data_mid_68_imag <= _zz_6221[15 : 0];
        data_mid_64_real <= _zz_6225[15 : 0];
        data_mid_64_imag <= _zz_6229[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_69_real <= _zz_6239[15 : 0];
        data_mid_69_imag <= _zz_6243[15 : 0];
        data_mid_65_real <= _zz_6247[15 : 0];
        data_mid_65_imag <= _zz_6251[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_70_real <= _zz_6261[15 : 0];
        data_mid_70_imag <= _zz_6265[15 : 0];
        data_mid_66_real <= _zz_6269[15 : 0];
        data_mid_66_imag <= _zz_6273[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_71_real <= _zz_6283[15 : 0];
        data_mid_71_imag <= _zz_6287[15 : 0];
        data_mid_67_real <= _zz_6291[15 : 0];
        data_mid_67_imag <= _zz_6295[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_76_real <= _zz_6305[15 : 0];
        data_mid_76_imag <= _zz_6309[15 : 0];
        data_mid_72_real <= _zz_6313[15 : 0];
        data_mid_72_imag <= _zz_6317[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_77_real <= _zz_6327[15 : 0];
        data_mid_77_imag <= _zz_6331[15 : 0];
        data_mid_73_real <= _zz_6335[15 : 0];
        data_mid_73_imag <= _zz_6339[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_78_real <= _zz_6349[15 : 0];
        data_mid_78_imag <= _zz_6353[15 : 0];
        data_mid_74_real <= _zz_6357[15 : 0];
        data_mid_74_imag <= _zz_6361[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_79_real <= _zz_6371[15 : 0];
        data_mid_79_imag <= _zz_6375[15 : 0];
        data_mid_75_real <= _zz_6379[15 : 0];
        data_mid_75_imag <= _zz_6383[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_84_real <= _zz_6393[15 : 0];
        data_mid_84_imag <= _zz_6397[15 : 0];
        data_mid_80_real <= _zz_6401[15 : 0];
        data_mid_80_imag <= _zz_6405[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_85_real <= _zz_6415[15 : 0];
        data_mid_85_imag <= _zz_6419[15 : 0];
        data_mid_81_real <= _zz_6423[15 : 0];
        data_mid_81_imag <= _zz_6427[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_86_real <= _zz_6437[15 : 0];
        data_mid_86_imag <= _zz_6441[15 : 0];
        data_mid_82_real <= _zz_6445[15 : 0];
        data_mid_82_imag <= _zz_6449[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_87_real <= _zz_6459[15 : 0];
        data_mid_87_imag <= _zz_6463[15 : 0];
        data_mid_83_real <= _zz_6467[15 : 0];
        data_mid_83_imag <= _zz_6471[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_92_real <= _zz_6481[15 : 0];
        data_mid_92_imag <= _zz_6485[15 : 0];
        data_mid_88_real <= _zz_6489[15 : 0];
        data_mid_88_imag <= _zz_6493[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_93_real <= _zz_6503[15 : 0];
        data_mid_93_imag <= _zz_6507[15 : 0];
        data_mid_89_real <= _zz_6511[15 : 0];
        data_mid_89_imag <= _zz_6515[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_94_real <= _zz_6525[15 : 0];
        data_mid_94_imag <= _zz_6529[15 : 0];
        data_mid_90_real <= _zz_6533[15 : 0];
        data_mid_90_imag <= _zz_6537[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_95_real <= _zz_6547[15 : 0];
        data_mid_95_imag <= _zz_6551[15 : 0];
        data_mid_91_real <= _zz_6555[15 : 0];
        data_mid_91_imag <= _zz_6559[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_100_real <= _zz_6569[15 : 0];
        data_mid_100_imag <= _zz_6573[15 : 0];
        data_mid_96_real <= _zz_6577[15 : 0];
        data_mid_96_imag <= _zz_6581[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_101_real <= _zz_6591[15 : 0];
        data_mid_101_imag <= _zz_6595[15 : 0];
        data_mid_97_real <= _zz_6599[15 : 0];
        data_mid_97_imag <= _zz_6603[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_102_real <= _zz_6613[15 : 0];
        data_mid_102_imag <= _zz_6617[15 : 0];
        data_mid_98_real <= _zz_6621[15 : 0];
        data_mid_98_imag <= _zz_6625[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_103_real <= _zz_6635[15 : 0];
        data_mid_103_imag <= _zz_6639[15 : 0];
        data_mid_99_real <= _zz_6643[15 : 0];
        data_mid_99_imag <= _zz_6647[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_108_real <= _zz_6657[15 : 0];
        data_mid_108_imag <= _zz_6661[15 : 0];
        data_mid_104_real <= _zz_6665[15 : 0];
        data_mid_104_imag <= _zz_6669[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_109_real <= _zz_6679[15 : 0];
        data_mid_109_imag <= _zz_6683[15 : 0];
        data_mid_105_real <= _zz_6687[15 : 0];
        data_mid_105_imag <= _zz_6691[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_110_real <= _zz_6701[15 : 0];
        data_mid_110_imag <= _zz_6705[15 : 0];
        data_mid_106_real <= _zz_6709[15 : 0];
        data_mid_106_imag <= _zz_6713[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_111_real <= _zz_6723[15 : 0];
        data_mid_111_imag <= _zz_6727[15 : 0];
        data_mid_107_real <= _zz_6731[15 : 0];
        data_mid_107_imag <= _zz_6735[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_116_real <= _zz_6745[15 : 0];
        data_mid_116_imag <= _zz_6749[15 : 0];
        data_mid_112_real <= _zz_6753[15 : 0];
        data_mid_112_imag <= _zz_6757[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_117_real <= _zz_6767[15 : 0];
        data_mid_117_imag <= _zz_6771[15 : 0];
        data_mid_113_real <= _zz_6775[15 : 0];
        data_mid_113_imag <= _zz_6779[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_118_real <= _zz_6789[15 : 0];
        data_mid_118_imag <= _zz_6793[15 : 0];
        data_mid_114_real <= _zz_6797[15 : 0];
        data_mid_114_imag <= _zz_6801[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_119_real <= _zz_6811[15 : 0];
        data_mid_119_imag <= _zz_6815[15 : 0];
        data_mid_115_real <= _zz_6819[15 : 0];
        data_mid_115_imag <= _zz_6823[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_124_real <= _zz_6833[15 : 0];
        data_mid_124_imag <= _zz_6837[15 : 0];
        data_mid_120_real <= _zz_6841[15 : 0];
        data_mid_120_imag <= _zz_6845[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_125_real <= _zz_6855[15 : 0];
        data_mid_125_imag <= _zz_6859[15 : 0];
        data_mid_121_real <= _zz_6863[15 : 0];
        data_mid_121_imag <= _zz_6867[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_126_real <= _zz_6877[15 : 0];
        data_mid_126_imag <= _zz_6881[15 : 0];
        data_mid_122_real <= _zz_6885[15 : 0];
        data_mid_122_imag <= _zz_6889[15 : 0];
      end
      if((current_level_cnt_value == 3'b011))begin
        data_mid_127_real <= _zz_6899[15 : 0];
        data_mid_127_imag <= _zz_6903[15 : 0];
        data_mid_123_real <= _zz_6907[15 : 0];
        data_mid_123_imag <= _zz_6911[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_8_real <= _zz_6921[15 : 0];
        data_mid_8_imag <= _zz_6925[15 : 0];
        data_mid_0_real <= _zz_6929[15 : 0];
        data_mid_0_imag <= _zz_6933[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_9_real <= _zz_6943[15 : 0];
        data_mid_9_imag <= _zz_6947[15 : 0];
        data_mid_1_real <= _zz_6951[15 : 0];
        data_mid_1_imag <= _zz_6955[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_10_real <= _zz_6965[15 : 0];
        data_mid_10_imag <= _zz_6969[15 : 0];
        data_mid_2_real <= _zz_6973[15 : 0];
        data_mid_2_imag <= _zz_6977[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_11_real <= _zz_6987[15 : 0];
        data_mid_11_imag <= _zz_6991[15 : 0];
        data_mid_3_real <= _zz_6995[15 : 0];
        data_mid_3_imag <= _zz_6999[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_12_real <= _zz_7009[15 : 0];
        data_mid_12_imag <= _zz_7013[15 : 0];
        data_mid_4_real <= _zz_7017[15 : 0];
        data_mid_4_imag <= _zz_7021[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_13_real <= _zz_7031[15 : 0];
        data_mid_13_imag <= _zz_7035[15 : 0];
        data_mid_5_real <= _zz_7039[15 : 0];
        data_mid_5_imag <= _zz_7043[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_14_real <= _zz_7053[15 : 0];
        data_mid_14_imag <= _zz_7057[15 : 0];
        data_mid_6_real <= _zz_7061[15 : 0];
        data_mid_6_imag <= _zz_7065[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_15_real <= _zz_7075[15 : 0];
        data_mid_15_imag <= _zz_7079[15 : 0];
        data_mid_7_real <= _zz_7083[15 : 0];
        data_mid_7_imag <= _zz_7087[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_24_real <= _zz_7097[15 : 0];
        data_mid_24_imag <= _zz_7101[15 : 0];
        data_mid_16_real <= _zz_7105[15 : 0];
        data_mid_16_imag <= _zz_7109[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_25_real <= _zz_7119[15 : 0];
        data_mid_25_imag <= _zz_7123[15 : 0];
        data_mid_17_real <= _zz_7127[15 : 0];
        data_mid_17_imag <= _zz_7131[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_26_real <= _zz_7141[15 : 0];
        data_mid_26_imag <= _zz_7145[15 : 0];
        data_mid_18_real <= _zz_7149[15 : 0];
        data_mid_18_imag <= _zz_7153[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_27_real <= _zz_7163[15 : 0];
        data_mid_27_imag <= _zz_7167[15 : 0];
        data_mid_19_real <= _zz_7171[15 : 0];
        data_mid_19_imag <= _zz_7175[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_28_real <= _zz_7185[15 : 0];
        data_mid_28_imag <= _zz_7189[15 : 0];
        data_mid_20_real <= _zz_7193[15 : 0];
        data_mid_20_imag <= _zz_7197[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_29_real <= _zz_7207[15 : 0];
        data_mid_29_imag <= _zz_7211[15 : 0];
        data_mid_21_real <= _zz_7215[15 : 0];
        data_mid_21_imag <= _zz_7219[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_30_real <= _zz_7229[15 : 0];
        data_mid_30_imag <= _zz_7233[15 : 0];
        data_mid_22_real <= _zz_7237[15 : 0];
        data_mid_22_imag <= _zz_7241[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_31_real <= _zz_7251[15 : 0];
        data_mid_31_imag <= _zz_7255[15 : 0];
        data_mid_23_real <= _zz_7259[15 : 0];
        data_mid_23_imag <= _zz_7263[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_40_real <= _zz_7273[15 : 0];
        data_mid_40_imag <= _zz_7277[15 : 0];
        data_mid_32_real <= _zz_7281[15 : 0];
        data_mid_32_imag <= _zz_7285[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_41_real <= _zz_7295[15 : 0];
        data_mid_41_imag <= _zz_7299[15 : 0];
        data_mid_33_real <= _zz_7303[15 : 0];
        data_mid_33_imag <= _zz_7307[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_42_real <= _zz_7317[15 : 0];
        data_mid_42_imag <= _zz_7321[15 : 0];
        data_mid_34_real <= _zz_7325[15 : 0];
        data_mid_34_imag <= _zz_7329[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_43_real <= _zz_7339[15 : 0];
        data_mid_43_imag <= _zz_7343[15 : 0];
        data_mid_35_real <= _zz_7347[15 : 0];
        data_mid_35_imag <= _zz_7351[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_44_real <= _zz_7361[15 : 0];
        data_mid_44_imag <= _zz_7365[15 : 0];
        data_mid_36_real <= _zz_7369[15 : 0];
        data_mid_36_imag <= _zz_7373[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_45_real <= _zz_7383[15 : 0];
        data_mid_45_imag <= _zz_7387[15 : 0];
        data_mid_37_real <= _zz_7391[15 : 0];
        data_mid_37_imag <= _zz_7395[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_46_real <= _zz_7405[15 : 0];
        data_mid_46_imag <= _zz_7409[15 : 0];
        data_mid_38_real <= _zz_7413[15 : 0];
        data_mid_38_imag <= _zz_7417[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_47_real <= _zz_7427[15 : 0];
        data_mid_47_imag <= _zz_7431[15 : 0];
        data_mid_39_real <= _zz_7435[15 : 0];
        data_mid_39_imag <= _zz_7439[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_56_real <= _zz_7449[15 : 0];
        data_mid_56_imag <= _zz_7453[15 : 0];
        data_mid_48_real <= _zz_7457[15 : 0];
        data_mid_48_imag <= _zz_7461[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_57_real <= _zz_7471[15 : 0];
        data_mid_57_imag <= _zz_7475[15 : 0];
        data_mid_49_real <= _zz_7479[15 : 0];
        data_mid_49_imag <= _zz_7483[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_58_real <= _zz_7493[15 : 0];
        data_mid_58_imag <= _zz_7497[15 : 0];
        data_mid_50_real <= _zz_7501[15 : 0];
        data_mid_50_imag <= _zz_7505[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_59_real <= _zz_7515[15 : 0];
        data_mid_59_imag <= _zz_7519[15 : 0];
        data_mid_51_real <= _zz_7523[15 : 0];
        data_mid_51_imag <= _zz_7527[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_60_real <= _zz_7537[15 : 0];
        data_mid_60_imag <= _zz_7541[15 : 0];
        data_mid_52_real <= _zz_7545[15 : 0];
        data_mid_52_imag <= _zz_7549[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_61_real <= _zz_7559[15 : 0];
        data_mid_61_imag <= _zz_7563[15 : 0];
        data_mid_53_real <= _zz_7567[15 : 0];
        data_mid_53_imag <= _zz_7571[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_62_real <= _zz_7581[15 : 0];
        data_mid_62_imag <= _zz_7585[15 : 0];
        data_mid_54_real <= _zz_7589[15 : 0];
        data_mid_54_imag <= _zz_7593[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_63_real <= _zz_7603[15 : 0];
        data_mid_63_imag <= _zz_7607[15 : 0];
        data_mid_55_real <= _zz_7611[15 : 0];
        data_mid_55_imag <= _zz_7615[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_72_real <= _zz_7625[15 : 0];
        data_mid_72_imag <= _zz_7629[15 : 0];
        data_mid_64_real <= _zz_7633[15 : 0];
        data_mid_64_imag <= _zz_7637[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_73_real <= _zz_7647[15 : 0];
        data_mid_73_imag <= _zz_7651[15 : 0];
        data_mid_65_real <= _zz_7655[15 : 0];
        data_mid_65_imag <= _zz_7659[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_74_real <= _zz_7669[15 : 0];
        data_mid_74_imag <= _zz_7673[15 : 0];
        data_mid_66_real <= _zz_7677[15 : 0];
        data_mid_66_imag <= _zz_7681[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_75_real <= _zz_7691[15 : 0];
        data_mid_75_imag <= _zz_7695[15 : 0];
        data_mid_67_real <= _zz_7699[15 : 0];
        data_mid_67_imag <= _zz_7703[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_76_real <= _zz_7713[15 : 0];
        data_mid_76_imag <= _zz_7717[15 : 0];
        data_mid_68_real <= _zz_7721[15 : 0];
        data_mid_68_imag <= _zz_7725[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_77_real <= _zz_7735[15 : 0];
        data_mid_77_imag <= _zz_7739[15 : 0];
        data_mid_69_real <= _zz_7743[15 : 0];
        data_mid_69_imag <= _zz_7747[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_78_real <= _zz_7757[15 : 0];
        data_mid_78_imag <= _zz_7761[15 : 0];
        data_mid_70_real <= _zz_7765[15 : 0];
        data_mid_70_imag <= _zz_7769[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_79_real <= _zz_7779[15 : 0];
        data_mid_79_imag <= _zz_7783[15 : 0];
        data_mid_71_real <= _zz_7787[15 : 0];
        data_mid_71_imag <= _zz_7791[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_88_real <= _zz_7801[15 : 0];
        data_mid_88_imag <= _zz_7805[15 : 0];
        data_mid_80_real <= _zz_7809[15 : 0];
        data_mid_80_imag <= _zz_7813[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_89_real <= _zz_7823[15 : 0];
        data_mid_89_imag <= _zz_7827[15 : 0];
        data_mid_81_real <= _zz_7831[15 : 0];
        data_mid_81_imag <= _zz_7835[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_90_real <= _zz_7845[15 : 0];
        data_mid_90_imag <= _zz_7849[15 : 0];
        data_mid_82_real <= _zz_7853[15 : 0];
        data_mid_82_imag <= _zz_7857[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_91_real <= _zz_7867[15 : 0];
        data_mid_91_imag <= _zz_7871[15 : 0];
        data_mid_83_real <= _zz_7875[15 : 0];
        data_mid_83_imag <= _zz_7879[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_92_real <= _zz_7889[15 : 0];
        data_mid_92_imag <= _zz_7893[15 : 0];
        data_mid_84_real <= _zz_7897[15 : 0];
        data_mid_84_imag <= _zz_7901[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_93_real <= _zz_7911[15 : 0];
        data_mid_93_imag <= _zz_7915[15 : 0];
        data_mid_85_real <= _zz_7919[15 : 0];
        data_mid_85_imag <= _zz_7923[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_94_real <= _zz_7933[15 : 0];
        data_mid_94_imag <= _zz_7937[15 : 0];
        data_mid_86_real <= _zz_7941[15 : 0];
        data_mid_86_imag <= _zz_7945[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_95_real <= _zz_7955[15 : 0];
        data_mid_95_imag <= _zz_7959[15 : 0];
        data_mid_87_real <= _zz_7963[15 : 0];
        data_mid_87_imag <= _zz_7967[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_104_real <= _zz_7977[15 : 0];
        data_mid_104_imag <= _zz_7981[15 : 0];
        data_mid_96_real <= _zz_7985[15 : 0];
        data_mid_96_imag <= _zz_7989[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_105_real <= _zz_7999[15 : 0];
        data_mid_105_imag <= _zz_8003[15 : 0];
        data_mid_97_real <= _zz_8007[15 : 0];
        data_mid_97_imag <= _zz_8011[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_106_real <= _zz_8021[15 : 0];
        data_mid_106_imag <= _zz_8025[15 : 0];
        data_mid_98_real <= _zz_8029[15 : 0];
        data_mid_98_imag <= _zz_8033[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_107_real <= _zz_8043[15 : 0];
        data_mid_107_imag <= _zz_8047[15 : 0];
        data_mid_99_real <= _zz_8051[15 : 0];
        data_mid_99_imag <= _zz_8055[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_108_real <= _zz_8065[15 : 0];
        data_mid_108_imag <= _zz_8069[15 : 0];
        data_mid_100_real <= _zz_8073[15 : 0];
        data_mid_100_imag <= _zz_8077[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_109_real <= _zz_8087[15 : 0];
        data_mid_109_imag <= _zz_8091[15 : 0];
        data_mid_101_real <= _zz_8095[15 : 0];
        data_mid_101_imag <= _zz_8099[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_110_real <= _zz_8109[15 : 0];
        data_mid_110_imag <= _zz_8113[15 : 0];
        data_mid_102_real <= _zz_8117[15 : 0];
        data_mid_102_imag <= _zz_8121[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_111_real <= _zz_8131[15 : 0];
        data_mid_111_imag <= _zz_8135[15 : 0];
        data_mid_103_real <= _zz_8139[15 : 0];
        data_mid_103_imag <= _zz_8143[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_120_real <= _zz_8153[15 : 0];
        data_mid_120_imag <= _zz_8157[15 : 0];
        data_mid_112_real <= _zz_8161[15 : 0];
        data_mid_112_imag <= _zz_8165[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_121_real <= _zz_8175[15 : 0];
        data_mid_121_imag <= _zz_8179[15 : 0];
        data_mid_113_real <= _zz_8183[15 : 0];
        data_mid_113_imag <= _zz_8187[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_122_real <= _zz_8197[15 : 0];
        data_mid_122_imag <= _zz_8201[15 : 0];
        data_mid_114_real <= _zz_8205[15 : 0];
        data_mid_114_imag <= _zz_8209[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_123_real <= _zz_8219[15 : 0];
        data_mid_123_imag <= _zz_8223[15 : 0];
        data_mid_115_real <= _zz_8227[15 : 0];
        data_mid_115_imag <= _zz_8231[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_124_real <= _zz_8241[15 : 0];
        data_mid_124_imag <= _zz_8245[15 : 0];
        data_mid_116_real <= _zz_8249[15 : 0];
        data_mid_116_imag <= _zz_8253[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_125_real <= _zz_8263[15 : 0];
        data_mid_125_imag <= _zz_8267[15 : 0];
        data_mid_117_real <= _zz_8271[15 : 0];
        data_mid_117_imag <= _zz_8275[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_126_real <= _zz_8285[15 : 0];
        data_mid_126_imag <= _zz_8289[15 : 0];
        data_mid_118_real <= _zz_8293[15 : 0];
        data_mid_118_imag <= _zz_8297[15 : 0];
      end
      if((current_level_cnt_value == 3'b100))begin
        data_mid_127_real <= _zz_8307[15 : 0];
        data_mid_127_imag <= _zz_8311[15 : 0];
        data_mid_119_real <= _zz_8315[15 : 0];
        data_mid_119_imag <= _zz_8319[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_16_real <= _zz_8329[15 : 0];
        data_mid_16_imag <= _zz_8333[15 : 0];
        data_mid_0_real <= _zz_8337[15 : 0];
        data_mid_0_imag <= _zz_8341[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_17_real <= _zz_8351[15 : 0];
        data_mid_17_imag <= _zz_8355[15 : 0];
        data_mid_1_real <= _zz_8359[15 : 0];
        data_mid_1_imag <= _zz_8363[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_18_real <= _zz_8373[15 : 0];
        data_mid_18_imag <= _zz_8377[15 : 0];
        data_mid_2_real <= _zz_8381[15 : 0];
        data_mid_2_imag <= _zz_8385[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_19_real <= _zz_8395[15 : 0];
        data_mid_19_imag <= _zz_8399[15 : 0];
        data_mid_3_real <= _zz_8403[15 : 0];
        data_mid_3_imag <= _zz_8407[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_20_real <= _zz_8417[15 : 0];
        data_mid_20_imag <= _zz_8421[15 : 0];
        data_mid_4_real <= _zz_8425[15 : 0];
        data_mid_4_imag <= _zz_8429[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_21_real <= _zz_8439[15 : 0];
        data_mid_21_imag <= _zz_8443[15 : 0];
        data_mid_5_real <= _zz_8447[15 : 0];
        data_mid_5_imag <= _zz_8451[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_22_real <= _zz_8461[15 : 0];
        data_mid_22_imag <= _zz_8465[15 : 0];
        data_mid_6_real <= _zz_8469[15 : 0];
        data_mid_6_imag <= _zz_8473[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_23_real <= _zz_8483[15 : 0];
        data_mid_23_imag <= _zz_8487[15 : 0];
        data_mid_7_real <= _zz_8491[15 : 0];
        data_mid_7_imag <= _zz_8495[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_24_real <= _zz_8505[15 : 0];
        data_mid_24_imag <= _zz_8509[15 : 0];
        data_mid_8_real <= _zz_8513[15 : 0];
        data_mid_8_imag <= _zz_8517[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_25_real <= _zz_8527[15 : 0];
        data_mid_25_imag <= _zz_8531[15 : 0];
        data_mid_9_real <= _zz_8535[15 : 0];
        data_mid_9_imag <= _zz_8539[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_26_real <= _zz_8549[15 : 0];
        data_mid_26_imag <= _zz_8553[15 : 0];
        data_mid_10_real <= _zz_8557[15 : 0];
        data_mid_10_imag <= _zz_8561[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_27_real <= _zz_8571[15 : 0];
        data_mid_27_imag <= _zz_8575[15 : 0];
        data_mid_11_real <= _zz_8579[15 : 0];
        data_mid_11_imag <= _zz_8583[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_28_real <= _zz_8593[15 : 0];
        data_mid_28_imag <= _zz_8597[15 : 0];
        data_mid_12_real <= _zz_8601[15 : 0];
        data_mid_12_imag <= _zz_8605[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_29_real <= _zz_8615[15 : 0];
        data_mid_29_imag <= _zz_8619[15 : 0];
        data_mid_13_real <= _zz_8623[15 : 0];
        data_mid_13_imag <= _zz_8627[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_30_real <= _zz_8637[15 : 0];
        data_mid_30_imag <= _zz_8641[15 : 0];
        data_mid_14_real <= _zz_8645[15 : 0];
        data_mid_14_imag <= _zz_8649[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_31_real <= _zz_8659[15 : 0];
        data_mid_31_imag <= _zz_8663[15 : 0];
        data_mid_15_real <= _zz_8667[15 : 0];
        data_mid_15_imag <= _zz_8671[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_48_real <= _zz_8681[15 : 0];
        data_mid_48_imag <= _zz_8685[15 : 0];
        data_mid_32_real <= _zz_8689[15 : 0];
        data_mid_32_imag <= _zz_8693[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_49_real <= _zz_8703[15 : 0];
        data_mid_49_imag <= _zz_8707[15 : 0];
        data_mid_33_real <= _zz_8711[15 : 0];
        data_mid_33_imag <= _zz_8715[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_50_real <= _zz_8725[15 : 0];
        data_mid_50_imag <= _zz_8729[15 : 0];
        data_mid_34_real <= _zz_8733[15 : 0];
        data_mid_34_imag <= _zz_8737[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_51_real <= _zz_8747[15 : 0];
        data_mid_51_imag <= _zz_8751[15 : 0];
        data_mid_35_real <= _zz_8755[15 : 0];
        data_mid_35_imag <= _zz_8759[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_52_real <= _zz_8769[15 : 0];
        data_mid_52_imag <= _zz_8773[15 : 0];
        data_mid_36_real <= _zz_8777[15 : 0];
        data_mid_36_imag <= _zz_8781[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_53_real <= _zz_8791[15 : 0];
        data_mid_53_imag <= _zz_8795[15 : 0];
        data_mid_37_real <= _zz_8799[15 : 0];
        data_mid_37_imag <= _zz_8803[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_54_real <= _zz_8813[15 : 0];
        data_mid_54_imag <= _zz_8817[15 : 0];
        data_mid_38_real <= _zz_8821[15 : 0];
        data_mid_38_imag <= _zz_8825[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_55_real <= _zz_8835[15 : 0];
        data_mid_55_imag <= _zz_8839[15 : 0];
        data_mid_39_real <= _zz_8843[15 : 0];
        data_mid_39_imag <= _zz_8847[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_56_real <= _zz_8857[15 : 0];
        data_mid_56_imag <= _zz_8861[15 : 0];
        data_mid_40_real <= _zz_8865[15 : 0];
        data_mid_40_imag <= _zz_8869[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_57_real <= _zz_8879[15 : 0];
        data_mid_57_imag <= _zz_8883[15 : 0];
        data_mid_41_real <= _zz_8887[15 : 0];
        data_mid_41_imag <= _zz_8891[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_58_real <= _zz_8901[15 : 0];
        data_mid_58_imag <= _zz_8905[15 : 0];
        data_mid_42_real <= _zz_8909[15 : 0];
        data_mid_42_imag <= _zz_8913[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_59_real <= _zz_8923[15 : 0];
        data_mid_59_imag <= _zz_8927[15 : 0];
        data_mid_43_real <= _zz_8931[15 : 0];
        data_mid_43_imag <= _zz_8935[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_60_real <= _zz_8945[15 : 0];
        data_mid_60_imag <= _zz_8949[15 : 0];
        data_mid_44_real <= _zz_8953[15 : 0];
        data_mid_44_imag <= _zz_8957[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_61_real <= _zz_8967[15 : 0];
        data_mid_61_imag <= _zz_8971[15 : 0];
        data_mid_45_real <= _zz_8975[15 : 0];
        data_mid_45_imag <= _zz_8979[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_62_real <= _zz_8989[15 : 0];
        data_mid_62_imag <= _zz_8993[15 : 0];
        data_mid_46_real <= _zz_8997[15 : 0];
        data_mid_46_imag <= _zz_9001[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_63_real <= _zz_9011[15 : 0];
        data_mid_63_imag <= _zz_9015[15 : 0];
        data_mid_47_real <= _zz_9019[15 : 0];
        data_mid_47_imag <= _zz_9023[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_80_real <= _zz_9033[15 : 0];
        data_mid_80_imag <= _zz_9037[15 : 0];
        data_mid_64_real <= _zz_9041[15 : 0];
        data_mid_64_imag <= _zz_9045[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_81_real <= _zz_9055[15 : 0];
        data_mid_81_imag <= _zz_9059[15 : 0];
        data_mid_65_real <= _zz_9063[15 : 0];
        data_mid_65_imag <= _zz_9067[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_82_real <= _zz_9077[15 : 0];
        data_mid_82_imag <= _zz_9081[15 : 0];
        data_mid_66_real <= _zz_9085[15 : 0];
        data_mid_66_imag <= _zz_9089[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_83_real <= _zz_9099[15 : 0];
        data_mid_83_imag <= _zz_9103[15 : 0];
        data_mid_67_real <= _zz_9107[15 : 0];
        data_mid_67_imag <= _zz_9111[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_84_real <= _zz_9121[15 : 0];
        data_mid_84_imag <= _zz_9125[15 : 0];
        data_mid_68_real <= _zz_9129[15 : 0];
        data_mid_68_imag <= _zz_9133[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_85_real <= _zz_9143[15 : 0];
        data_mid_85_imag <= _zz_9147[15 : 0];
        data_mid_69_real <= _zz_9151[15 : 0];
        data_mid_69_imag <= _zz_9155[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_86_real <= _zz_9165[15 : 0];
        data_mid_86_imag <= _zz_9169[15 : 0];
        data_mid_70_real <= _zz_9173[15 : 0];
        data_mid_70_imag <= _zz_9177[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_87_real <= _zz_9187[15 : 0];
        data_mid_87_imag <= _zz_9191[15 : 0];
        data_mid_71_real <= _zz_9195[15 : 0];
        data_mid_71_imag <= _zz_9199[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_88_real <= _zz_9209[15 : 0];
        data_mid_88_imag <= _zz_9213[15 : 0];
        data_mid_72_real <= _zz_9217[15 : 0];
        data_mid_72_imag <= _zz_9221[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_89_real <= _zz_9231[15 : 0];
        data_mid_89_imag <= _zz_9235[15 : 0];
        data_mid_73_real <= _zz_9239[15 : 0];
        data_mid_73_imag <= _zz_9243[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_90_real <= _zz_9253[15 : 0];
        data_mid_90_imag <= _zz_9257[15 : 0];
        data_mid_74_real <= _zz_9261[15 : 0];
        data_mid_74_imag <= _zz_9265[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_91_real <= _zz_9275[15 : 0];
        data_mid_91_imag <= _zz_9279[15 : 0];
        data_mid_75_real <= _zz_9283[15 : 0];
        data_mid_75_imag <= _zz_9287[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_92_real <= _zz_9297[15 : 0];
        data_mid_92_imag <= _zz_9301[15 : 0];
        data_mid_76_real <= _zz_9305[15 : 0];
        data_mid_76_imag <= _zz_9309[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_93_real <= _zz_9319[15 : 0];
        data_mid_93_imag <= _zz_9323[15 : 0];
        data_mid_77_real <= _zz_9327[15 : 0];
        data_mid_77_imag <= _zz_9331[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_94_real <= _zz_9341[15 : 0];
        data_mid_94_imag <= _zz_9345[15 : 0];
        data_mid_78_real <= _zz_9349[15 : 0];
        data_mid_78_imag <= _zz_9353[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_95_real <= _zz_9363[15 : 0];
        data_mid_95_imag <= _zz_9367[15 : 0];
        data_mid_79_real <= _zz_9371[15 : 0];
        data_mid_79_imag <= _zz_9375[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_112_real <= _zz_9385[15 : 0];
        data_mid_112_imag <= _zz_9389[15 : 0];
        data_mid_96_real <= _zz_9393[15 : 0];
        data_mid_96_imag <= _zz_9397[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_113_real <= _zz_9407[15 : 0];
        data_mid_113_imag <= _zz_9411[15 : 0];
        data_mid_97_real <= _zz_9415[15 : 0];
        data_mid_97_imag <= _zz_9419[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_114_real <= _zz_9429[15 : 0];
        data_mid_114_imag <= _zz_9433[15 : 0];
        data_mid_98_real <= _zz_9437[15 : 0];
        data_mid_98_imag <= _zz_9441[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_115_real <= _zz_9451[15 : 0];
        data_mid_115_imag <= _zz_9455[15 : 0];
        data_mid_99_real <= _zz_9459[15 : 0];
        data_mid_99_imag <= _zz_9463[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_116_real <= _zz_9473[15 : 0];
        data_mid_116_imag <= _zz_9477[15 : 0];
        data_mid_100_real <= _zz_9481[15 : 0];
        data_mid_100_imag <= _zz_9485[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_117_real <= _zz_9495[15 : 0];
        data_mid_117_imag <= _zz_9499[15 : 0];
        data_mid_101_real <= _zz_9503[15 : 0];
        data_mid_101_imag <= _zz_9507[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_118_real <= _zz_9517[15 : 0];
        data_mid_118_imag <= _zz_9521[15 : 0];
        data_mid_102_real <= _zz_9525[15 : 0];
        data_mid_102_imag <= _zz_9529[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_119_real <= _zz_9539[15 : 0];
        data_mid_119_imag <= _zz_9543[15 : 0];
        data_mid_103_real <= _zz_9547[15 : 0];
        data_mid_103_imag <= _zz_9551[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_120_real <= _zz_9561[15 : 0];
        data_mid_120_imag <= _zz_9565[15 : 0];
        data_mid_104_real <= _zz_9569[15 : 0];
        data_mid_104_imag <= _zz_9573[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_121_real <= _zz_9583[15 : 0];
        data_mid_121_imag <= _zz_9587[15 : 0];
        data_mid_105_real <= _zz_9591[15 : 0];
        data_mid_105_imag <= _zz_9595[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_122_real <= _zz_9605[15 : 0];
        data_mid_122_imag <= _zz_9609[15 : 0];
        data_mid_106_real <= _zz_9613[15 : 0];
        data_mid_106_imag <= _zz_9617[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_123_real <= _zz_9627[15 : 0];
        data_mid_123_imag <= _zz_9631[15 : 0];
        data_mid_107_real <= _zz_9635[15 : 0];
        data_mid_107_imag <= _zz_9639[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_124_real <= _zz_9649[15 : 0];
        data_mid_124_imag <= _zz_9653[15 : 0];
        data_mid_108_real <= _zz_9657[15 : 0];
        data_mid_108_imag <= _zz_9661[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_125_real <= _zz_9671[15 : 0];
        data_mid_125_imag <= _zz_9675[15 : 0];
        data_mid_109_real <= _zz_9679[15 : 0];
        data_mid_109_imag <= _zz_9683[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_126_real <= _zz_9693[15 : 0];
        data_mid_126_imag <= _zz_9697[15 : 0];
        data_mid_110_real <= _zz_9701[15 : 0];
        data_mid_110_imag <= _zz_9705[15 : 0];
      end
      if((current_level_cnt_value == 3'b101))begin
        data_mid_127_real <= _zz_9715[15 : 0];
        data_mid_127_imag <= _zz_9719[15 : 0];
        data_mid_111_real <= _zz_9723[15 : 0];
        data_mid_111_imag <= _zz_9727[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_32_real <= _zz_9737[15 : 0];
        data_mid_32_imag <= _zz_9741[15 : 0];
        data_mid_0_real <= _zz_9745[15 : 0];
        data_mid_0_imag <= _zz_9749[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_33_real <= _zz_9759[15 : 0];
        data_mid_33_imag <= _zz_9763[15 : 0];
        data_mid_1_real <= _zz_9767[15 : 0];
        data_mid_1_imag <= _zz_9771[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_34_real <= _zz_9781[15 : 0];
        data_mid_34_imag <= _zz_9785[15 : 0];
        data_mid_2_real <= _zz_9789[15 : 0];
        data_mid_2_imag <= _zz_9793[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_35_real <= _zz_9803[15 : 0];
        data_mid_35_imag <= _zz_9807[15 : 0];
        data_mid_3_real <= _zz_9811[15 : 0];
        data_mid_3_imag <= _zz_9815[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_36_real <= _zz_9825[15 : 0];
        data_mid_36_imag <= _zz_9829[15 : 0];
        data_mid_4_real <= _zz_9833[15 : 0];
        data_mid_4_imag <= _zz_9837[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_37_real <= _zz_9847[15 : 0];
        data_mid_37_imag <= _zz_9851[15 : 0];
        data_mid_5_real <= _zz_9855[15 : 0];
        data_mid_5_imag <= _zz_9859[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_38_real <= _zz_9869[15 : 0];
        data_mid_38_imag <= _zz_9873[15 : 0];
        data_mid_6_real <= _zz_9877[15 : 0];
        data_mid_6_imag <= _zz_9881[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_39_real <= _zz_9891[15 : 0];
        data_mid_39_imag <= _zz_9895[15 : 0];
        data_mid_7_real <= _zz_9899[15 : 0];
        data_mid_7_imag <= _zz_9903[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_40_real <= _zz_9913[15 : 0];
        data_mid_40_imag <= _zz_9917[15 : 0];
        data_mid_8_real <= _zz_9921[15 : 0];
        data_mid_8_imag <= _zz_9925[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_41_real <= _zz_9935[15 : 0];
        data_mid_41_imag <= _zz_9939[15 : 0];
        data_mid_9_real <= _zz_9943[15 : 0];
        data_mid_9_imag <= _zz_9947[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_42_real <= _zz_9957[15 : 0];
        data_mid_42_imag <= _zz_9961[15 : 0];
        data_mid_10_real <= _zz_9965[15 : 0];
        data_mid_10_imag <= _zz_9969[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_43_real <= _zz_9979[15 : 0];
        data_mid_43_imag <= _zz_9983[15 : 0];
        data_mid_11_real <= _zz_9987[15 : 0];
        data_mid_11_imag <= _zz_9991[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_44_real <= _zz_10001[15 : 0];
        data_mid_44_imag <= _zz_10005[15 : 0];
        data_mid_12_real <= _zz_10009[15 : 0];
        data_mid_12_imag <= _zz_10013[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_45_real <= _zz_10023[15 : 0];
        data_mid_45_imag <= _zz_10027[15 : 0];
        data_mid_13_real <= _zz_10031[15 : 0];
        data_mid_13_imag <= _zz_10035[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_46_real <= _zz_10045[15 : 0];
        data_mid_46_imag <= _zz_10049[15 : 0];
        data_mid_14_real <= _zz_10053[15 : 0];
        data_mid_14_imag <= _zz_10057[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_47_real <= _zz_10067[15 : 0];
        data_mid_47_imag <= _zz_10071[15 : 0];
        data_mid_15_real <= _zz_10075[15 : 0];
        data_mid_15_imag <= _zz_10079[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_48_real <= _zz_10089[15 : 0];
        data_mid_48_imag <= _zz_10093[15 : 0];
        data_mid_16_real <= _zz_10097[15 : 0];
        data_mid_16_imag <= _zz_10101[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_49_real <= _zz_10111[15 : 0];
        data_mid_49_imag <= _zz_10115[15 : 0];
        data_mid_17_real <= _zz_10119[15 : 0];
        data_mid_17_imag <= _zz_10123[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_50_real <= _zz_10133[15 : 0];
        data_mid_50_imag <= _zz_10137[15 : 0];
        data_mid_18_real <= _zz_10141[15 : 0];
        data_mid_18_imag <= _zz_10145[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_51_real <= _zz_10155[15 : 0];
        data_mid_51_imag <= _zz_10159[15 : 0];
        data_mid_19_real <= _zz_10163[15 : 0];
        data_mid_19_imag <= _zz_10167[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_52_real <= _zz_10177[15 : 0];
        data_mid_52_imag <= _zz_10181[15 : 0];
        data_mid_20_real <= _zz_10185[15 : 0];
        data_mid_20_imag <= _zz_10189[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_53_real <= _zz_10199[15 : 0];
        data_mid_53_imag <= _zz_10203[15 : 0];
        data_mid_21_real <= _zz_10207[15 : 0];
        data_mid_21_imag <= _zz_10211[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_54_real <= _zz_10221[15 : 0];
        data_mid_54_imag <= _zz_10225[15 : 0];
        data_mid_22_real <= _zz_10229[15 : 0];
        data_mid_22_imag <= _zz_10233[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_55_real <= _zz_10243[15 : 0];
        data_mid_55_imag <= _zz_10247[15 : 0];
        data_mid_23_real <= _zz_10251[15 : 0];
        data_mid_23_imag <= _zz_10255[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_56_real <= _zz_10265[15 : 0];
        data_mid_56_imag <= _zz_10269[15 : 0];
        data_mid_24_real <= _zz_10273[15 : 0];
        data_mid_24_imag <= _zz_10277[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_57_real <= _zz_10287[15 : 0];
        data_mid_57_imag <= _zz_10291[15 : 0];
        data_mid_25_real <= _zz_10295[15 : 0];
        data_mid_25_imag <= _zz_10299[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_58_real <= _zz_10309[15 : 0];
        data_mid_58_imag <= _zz_10313[15 : 0];
        data_mid_26_real <= _zz_10317[15 : 0];
        data_mid_26_imag <= _zz_10321[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_59_real <= _zz_10331[15 : 0];
        data_mid_59_imag <= _zz_10335[15 : 0];
        data_mid_27_real <= _zz_10339[15 : 0];
        data_mid_27_imag <= _zz_10343[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_60_real <= _zz_10353[15 : 0];
        data_mid_60_imag <= _zz_10357[15 : 0];
        data_mid_28_real <= _zz_10361[15 : 0];
        data_mid_28_imag <= _zz_10365[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_61_real <= _zz_10375[15 : 0];
        data_mid_61_imag <= _zz_10379[15 : 0];
        data_mid_29_real <= _zz_10383[15 : 0];
        data_mid_29_imag <= _zz_10387[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_62_real <= _zz_10397[15 : 0];
        data_mid_62_imag <= _zz_10401[15 : 0];
        data_mid_30_real <= _zz_10405[15 : 0];
        data_mid_30_imag <= _zz_10409[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_63_real <= _zz_10419[15 : 0];
        data_mid_63_imag <= _zz_10423[15 : 0];
        data_mid_31_real <= _zz_10427[15 : 0];
        data_mid_31_imag <= _zz_10431[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_96_real <= _zz_10441[15 : 0];
        data_mid_96_imag <= _zz_10445[15 : 0];
        data_mid_64_real <= _zz_10449[15 : 0];
        data_mid_64_imag <= _zz_10453[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_97_real <= _zz_10463[15 : 0];
        data_mid_97_imag <= _zz_10467[15 : 0];
        data_mid_65_real <= _zz_10471[15 : 0];
        data_mid_65_imag <= _zz_10475[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_98_real <= _zz_10485[15 : 0];
        data_mid_98_imag <= _zz_10489[15 : 0];
        data_mid_66_real <= _zz_10493[15 : 0];
        data_mid_66_imag <= _zz_10497[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_99_real <= _zz_10507[15 : 0];
        data_mid_99_imag <= _zz_10511[15 : 0];
        data_mid_67_real <= _zz_10515[15 : 0];
        data_mid_67_imag <= _zz_10519[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_100_real <= _zz_10529[15 : 0];
        data_mid_100_imag <= _zz_10533[15 : 0];
        data_mid_68_real <= _zz_10537[15 : 0];
        data_mid_68_imag <= _zz_10541[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_101_real <= _zz_10551[15 : 0];
        data_mid_101_imag <= _zz_10555[15 : 0];
        data_mid_69_real <= _zz_10559[15 : 0];
        data_mid_69_imag <= _zz_10563[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_102_real <= _zz_10573[15 : 0];
        data_mid_102_imag <= _zz_10577[15 : 0];
        data_mid_70_real <= _zz_10581[15 : 0];
        data_mid_70_imag <= _zz_10585[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_103_real <= _zz_10595[15 : 0];
        data_mid_103_imag <= _zz_10599[15 : 0];
        data_mid_71_real <= _zz_10603[15 : 0];
        data_mid_71_imag <= _zz_10607[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_104_real <= _zz_10617[15 : 0];
        data_mid_104_imag <= _zz_10621[15 : 0];
        data_mid_72_real <= _zz_10625[15 : 0];
        data_mid_72_imag <= _zz_10629[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_105_real <= _zz_10639[15 : 0];
        data_mid_105_imag <= _zz_10643[15 : 0];
        data_mid_73_real <= _zz_10647[15 : 0];
        data_mid_73_imag <= _zz_10651[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_106_real <= _zz_10661[15 : 0];
        data_mid_106_imag <= _zz_10665[15 : 0];
        data_mid_74_real <= _zz_10669[15 : 0];
        data_mid_74_imag <= _zz_10673[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_107_real <= _zz_10683[15 : 0];
        data_mid_107_imag <= _zz_10687[15 : 0];
        data_mid_75_real <= _zz_10691[15 : 0];
        data_mid_75_imag <= _zz_10695[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_108_real <= _zz_10705[15 : 0];
        data_mid_108_imag <= _zz_10709[15 : 0];
        data_mid_76_real <= _zz_10713[15 : 0];
        data_mid_76_imag <= _zz_10717[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_109_real <= _zz_10727[15 : 0];
        data_mid_109_imag <= _zz_10731[15 : 0];
        data_mid_77_real <= _zz_10735[15 : 0];
        data_mid_77_imag <= _zz_10739[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_110_real <= _zz_10749[15 : 0];
        data_mid_110_imag <= _zz_10753[15 : 0];
        data_mid_78_real <= _zz_10757[15 : 0];
        data_mid_78_imag <= _zz_10761[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_111_real <= _zz_10771[15 : 0];
        data_mid_111_imag <= _zz_10775[15 : 0];
        data_mid_79_real <= _zz_10779[15 : 0];
        data_mid_79_imag <= _zz_10783[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_112_real <= _zz_10793[15 : 0];
        data_mid_112_imag <= _zz_10797[15 : 0];
        data_mid_80_real <= _zz_10801[15 : 0];
        data_mid_80_imag <= _zz_10805[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_113_real <= _zz_10815[15 : 0];
        data_mid_113_imag <= _zz_10819[15 : 0];
        data_mid_81_real <= _zz_10823[15 : 0];
        data_mid_81_imag <= _zz_10827[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_114_real <= _zz_10837[15 : 0];
        data_mid_114_imag <= _zz_10841[15 : 0];
        data_mid_82_real <= _zz_10845[15 : 0];
        data_mid_82_imag <= _zz_10849[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_115_real <= _zz_10859[15 : 0];
        data_mid_115_imag <= _zz_10863[15 : 0];
        data_mid_83_real <= _zz_10867[15 : 0];
        data_mid_83_imag <= _zz_10871[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_116_real <= _zz_10881[15 : 0];
        data_mid_116_imag <= _zz_10885[15 : 0];
        data_mid_84_real <= _zz_10889[15 : 0];
        data_mid_84_imag <= _zz_10893[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_117_real <= _zz_10903[15 : 0];
        data_mid_117_imag <= _zz_10907[15 : 0];
        data_mid_85_real <= _zz_10911[15 : 0];
        data_mid_85_imag <= _zz_10915[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_118_real <= _zz_10925[15 : 0];
        data_mid_118_imag <= _zz_10929[15 : 0];
        data_mid_86_real <= _zz_10933[15 : 0];
        data_mid_86_imag <= _zz_10937[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_119_real <= _zz_10947[15 : 0];
        data_mid_119_imag <= _zz_10951[15 : 0];
        data_mid_87_real <= _zz_10955[15 : 0];
        data_mid_87_imag <= _zz_10959[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_120_real <= _zz_10969[15 : 0];
        data_mid_120_imag <= _zz_10973[15 : 0];
        data_mid_88_real <= _zz_10977[15 : 0];
        data_mid_88_imag <= _zz_10981[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_121_real <= _zz_10991[15 : 0];
        data_mid_121_imag <= _zz_10995[15 : 0];
        data_mid_89_real <= _zz_10999[15 : 0];
        data_mid_89_imag <= _zz_11003[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_122_real <= _zz_11013[15 : 0];
        data_mid_122_imag <= _zz_11017[15 : 0];
        data_mid_90_real <= _zz_11021[15 : 0];
        data_mid_90_imag <= _zz_11025[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_123_real <= _zz_11035[15 : 0];
        data_mid_123_imag <= _zz_11039[15 : 0];
        data_mid_91_real <= _zz_11043[15 : 0];
        data_mid_91_imag <= _zz_11047[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_124_real <= _zz_11057[15 : 0];
        data_mid_124_imag <= _zz_11061[15 : 0];
        data_mid_92_real <= _zz_11065[15 : 0];
        data_mid_92_imag <= _zz_11069[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_125_real <= _zz_11079[15 : 0];
        data_mid_125_imag <= _zz_11083[15 : 0];
        data_mid_93_real <= _zz_11087[15 : 0];
        data_mid_93_imag <= _zz_11091[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_126_real <= _zz_11101[15 : 0];
        data_mid_126_imag <= _zz_11105[15 : 0];
        data_mid_94_real <= _zz_11109[15 : 0];
        data_mid_94_imag <= _zz_11113[15 : 0];
      end
      if((current_level_cnt_value == 3'b110))begin
        data_mid_127_real <= _zz_11123[15 : 0];
        data_mid_127_imag <= _zz_11127[15 : 0];
        data_mid_95_real <= _zz_11131[15 : 0];
        data_mid_95_imag <= _zz_11135[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_64_real <= _zz_11145[15 : 0];
        data_mid_64_imag <= _zz_11149[15 : 0];
        data_mid_0_real <= _zz_11153[15 : 0];
        data_mid_0_imag <= _zz_11157[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_65_real <= _zz_11167[15 : 0];
        data_mid_65_imag <= _zz_11171[15 : 0];
        data_mid_1_real <= _zz_11175[15 : 0];
        data_mid_1_imag <= _zz_11179[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_66_real <= _zz_11189[15 : 0];
        data_mid_66_imag <= _zz_11193[15 : 0];
        data_mid_2_real <= _zz_11197[15 : 0];
        data_mid_2_imag <= _zz_11201[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_67_real <= _zz_11211[15 : 0];
        data_mid_67_imag <= _zz_11215[15 : 0];
        data_mid_3_real <= _zz_11219[15 : 0];
        data_mid_3_imag <= _zz_11223[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_68_real <= _zz_11233[15 : 0];
        data_mid_68_imag <= _zz_11237[15 : 0];
        data_mid_4_real <= _zz_11241[15 : 0];
        data_mid_4_imag <= _zz_11245[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_69_real <= _zz_11255[15 : 0];
        data_mid_69_imag <= _zz_11259[15 : 0];
        data_mid_5_real <= _zz_11263[15 : 0];
        data_mid_5_imag <= _zz_11267[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_70_real <= _zz_11277[15 : 0];
        data_mid_70_imag <= _zz_11281[15 : 0];
        data_mid_6_real <= _zz_11285[15 : 0];
        data_mid_6_imag <= _zz_11289[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_71_real <= _zz_11299[15 : 0];
        data_mid_71_imag <= _zz_11303[15 : 0];
        data_mid_7_real <= _zz_11307[15 : 0];
        data_mid_7_imag <= _zz_11311[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_72_real <= _zz_11321[15 : 0];
        data_mid_72_imag <= _zz_11325[15 : 0];
        data_mid_8_real <= _zz_11329[15 : 0];
        data_mid_8_imag <= _zz_11333[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_73_real <= _zz_11343[15 : 0];
        data_mid_73_imag <= _zz_11347[15 : 0];
        data_mid_9_real <= _zz_11351[15 : 0];
        data_mid_9_imag <= _zz_11355[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_74_real <= _zz_11365[15 : 0];
        data_mid_74_imag <= _zz_11369[15 : 0];
        data_mid_10_real <= _zz_11373[15 : 0];
        data_mid_10_imag <= _zz_11377[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_75_real <= _zz_11387[15 : 0];
        data_mid_75_imag <= _zz_11391[15 : 0];
        data_mid_11_real <= _zz_11395[15 : 0];
        data_mid_11_imag <= _zz_11399[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_76_real <= _zz_11409[15 : 0];
        data_mid_76_imag <= _zz_11413[15 : 0];
        data_mid_12_real <= _zz_11417[15 : 0];
        data_mid_12_imag <= _zz_11421[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_77_real <= _zz_11431[15 : 0];
        data_mid_77_imag <= _zz_11435[15 : 0];
        data_mid_13_real <= _zz_11439[15 : 0];
        data_mid_13_imag <= _zz_11443[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_78_real <= _zz_11453[15 : 0];
        data_mid_78_imag <= _zz_11457[15 : 0];
        data_mid_14_real <= _zz_11461[15 : 0];
        data_mid_14_imag <= _zz_11465[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_79_real <= _zz_11475[15 : 0];
        data_mid_79_imag <= _zz_11479[15 : 0];
        data_mid_15_real <= _zz_11483[15 : 0];
        data_mid_15_imag <= _zz_11487[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_80_real <= _zz_11497[15 : 0];
        data_mid_80_imag <= _zz_11501[15 : 0];
        data_mid_16_real <= _zz_11505[15 : 0];
        data_mid_16_imag <= _zz_11509[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_81_real <= _zz_11519[15 : 0];
        data_mid_81_imag <= _zz_11523[15 : 0];
        data_mid_17_real <= _zz_11527[15 : 0];
        data_mid_17_imag <= _zz_11531[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_82_real <= _zz_11541[15 : 0];
        data_mid_82_imag <= _zz_11545[15 : 0];
        data_mid_18_real <= _zz_11549[15 : 0];
        data_mid_18_imag <= _zz_11553[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_83_real <= _zz_11563[15 : 0];
        data_mid_83_imag <= _zz_11567[15 : 0];
        data_mid_19_real <= _zz_11571[15 : 0];
        data_mid_19_imag <= _zz_11575[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_84_real <= _zz_11585[15 : 0];
        data_mid_84_imag <= _zz_11589[15 : 0];
        data_mid_20_real <= _zz_11593[15 : 0];
        data_mid_20_imag <= _zz_11597[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_85_real <= _zz_11607[15 : 0];
        data_mid_85_imag <= _zz_11611[15 : 0];
        data_mid_21_real <= _zz_11615[15 : 0];
        data_mid_21_imag <= _zz_11619[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_86_real <= _zz_11629[15 : 0];
        data_mid_86_imag <= _zz_11633[15 : 0];
        data_mid_22_real <= _zz_11637[15 : 0];
        data_mid_22_imag <= _zz_11641[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_87_real <= _zz_11651[15 : 0];
        data_mid_87_imag <= _zz_11655[15 : 0];
        data_mid_23_real <= _zz_11659[15 : 0];
        data_mid_23_imag <= _zz_11663[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_88_real <= _zz_11673[15 : 0];
        data_mid_88_imag <= _zz_11677[15 : 0];
        data_mid_24_real <= _zz_11681[15 : 0];
        data_mid_24_imag <= _zz_11685[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_89_real <= _zz_11695[15 : 0];
        data_mid_89_imag <= _zz_11699[15 : 0];
        data_mid_25_real <= _zz_11703[15 : 0];
        data_mid_25_imag <= _zz_11707[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_90_real <= _zz_11717[15 : 0];
        data_mid_90_imag <= _zz_11721[15 : 0];
        data_mid_26_real <= _zz_11725[15 : 0];
        data_mid_26_imag <= _zz_11729[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_91_real <= _zz_11739[15 : 0];
        data_mid_91_imag <= _zz_11743[15 : 0];
        data_mid_27_real <= _zz_11747[15 : 0];
        data_mid_27_imag <= _zz_11751[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_92_real <= _zz_11761[15 : 0];
        data_mid_92_imag <= _zz_11765[15 : 0];
        data_mid_28_real <= _zz_11769[15 : 0];
        data_mid_28_imag <= _zz_11773[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_93_real <= _zz_11783[15 : 0];
        data_mid_93_imag <= _zz_11787[15 : 0];
        data_mid_29_real <= _zz_11791[15 : 0];
        data_mid_29_imag <= _zz_11795[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_94_real <= _zz_11805[15 : 0];
        data_mid_94_imag <= _zz_11809[15 : 0];
        data_mid_30_real <= _zz_11813[15 : 0];
        data_mid_30_imag <= _zz_11817[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_95_real <= _zz_11827[15 : 0];
        data_mid_95_imag <= _zz_11831[15 : 0];
        data_mid_31_real <= _zz_11835[15 : 0];
        data_mid_31_imag <= _zz_11839[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_96_real <= _zz_11849[15 : 0];
        data_mid_96_imag <= _zz_11853[15 : 0];
        data_mid_32_real <= _zz_11857[15 : 0];
        data_mid_32_imag <= _zz_11861[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_97_real <= _zz_11871[15 : 0];
        data_mid_97_imag <= _zz_11875[15 : 0];
        data_mid_33_real <= _zz_11879[15 : 0];
        data_mid_33_imag <= _zz_11883[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_98_real <= _zz_11893[15 : 0];
        data_mid_98_imag <= _zz_11897[15 : 0];
        data_mid_34_real <= _zz_11901[15 : 0];
        data_mid_34_imag <= _zz_11905[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_99_real <= _zz_11915[15 : 0];
        data_mid_99_imag <= _zz_11919[15 : 0];
        data_mid_35_real <= _zz_11923[15 : 0];
        data_mid_35_imag <= _zz_11927[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_100_real <= _zz_11937[15 : 0];
        data_mid_100_imag <= _zz_11941[15 : 0];
        data_mid_36_real <= _zz_11945[15 : 0];
        data_mid_36_imag <= _zz_11949[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_101_real <= _zz_11959[15 : 0];
        data_mid_101_imag <= _zz_11963[15 : 0];
        data_mid_37_real <= _zz_11967[15 : 0];
        data_mid_37_imag <= _zz_11971[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_102_real <= _zz_11981[15 : 0];
        data_mid_102_imag <= _zz_11985[15 : 0];
        data_mid_38_real <= _zz_11989[15 : 0];
        data_mid_38_imag <= _zz_11993[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_103_real <= _zz_12003[15 : 0];
        data_mid_103_imag <= _zz_12007[15 : 0];
        data_mid_39_real <= _zz_12011[15 : 0];
        data_mid_39_imag <= _zz_12015[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_104_real <= _zz_12025[15 : 0];
        data_mid_104_imag <= _zz_12029[15 : 0];
        data_mid_40_real <= _zz_12033[15 : 0];
        data_mid_40_imag <= _zz_12037[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_105_real <= _zz_12047[15 : 0];
        data_mid_105_imag <= _zz_12051[15 : 0];
        data_mid_41_real <= _zz_12055[15 : 0];
        data_mid_41_imag <= _zz_12059[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_106_real <= _zz_12069[15 : 0];
        data_mid_106_imag <= _zz_12073[15 : 0];
        data_mid_42_real <= _zz_12077[15 : 0];
        data_mid_42_imag <= _zz_12081[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_107_real <= _zz_12091[15 : 0];
        data_mid_107_imag <= _zz_12095[15 : 0];
        data_mid_43_real <= _zz_12099[15 : 0];
        data_mid_43_imag <= _zz_12103[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_108_real <= _zz_12113[15 : 0];
        data_mid_108_imag <= _zz_12117[15 : 0];
        data_mid_44_real <= _zz_12121[15 : 0];
        data_mid_44_imag <= _zz_12125[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_109_real <= _zz_12135[15 : 0];
        data_mid_109_imag <= _zz_12139[15 : 0];
        data_mid_45_real <= _zz_12143[15 : 0];
        data_mid_45_imag <= _zz_12147[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_110_real <= _zz_12157[15 : 0];
        data_mid_110_imag <= _zz_12161[15 : 0];
        data_mid_46_real <= _zz_12165[15 : 0];
        data_mid_46_imag <= _zz_12169[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_111_real <= _zz_12179[15 : 0];
        data_mid_111_imag <= _zz_12183[15 : 0];
        data_mid_47_real <= _zz_12187[15 : 0];
        data_mid_47_imag <= _zz_12191[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_112_real <= _zz_12201[15 : 0];
        data_mid_112_imag <= _zz_12205[15 : 0];
        data_mid_48_real <= _zz_12209[15 : 0];
        data_mid_48_imag <= _zz_12213[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_113_real <= _zz_12223[15 : 0];
        data_mid_113_imag <= _zz_12227[15 : 0];
        data_mid_49_real <= _zz_12231[15 : 0];
        data_mid_49_imag <= _zz_12235[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_114_real <= _zz_12245[15 : 0];
        data_mid_114_imag <= _zz_12249[15 : 0];
        data_mid_50_real <= _zz_12253[15 : 0];
        data_mid_50_imag <= _zz_12257[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_115_real <= _zz_12267[15 : 0];
        data_mid_115_imag <= _zz_12271[15 : 0];
        data_mid_51_real <= _zz_12275[15 : 0];
        data_mid_51_imag <= _zz_12279[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_116_real <= _zz_12289[15 : 0];
        data_mid_116_imag <= _zz_12293[15 : 0];
        data_mid_52_real <= _zz_12297[15 : 0];
        data_mid_52_imag <= _zz_12301[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_117_real <= _zz_12311[15 : 0];
        data_mid_117_imag <= _zz_12315[15 : 0];
        data_mid_53_real <= _zz_12319[15 : 0];
        data_mid_53_imag <= _zz_12323[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_118_real <= _zz_12333[15 : 0];
        data_mid_118_imag <= _zz_12337[15 : 0];
        data_mid_54_real <= _zz_12341[15 : 0];
        data_mid_54_imag <= _zz_12345[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_119_real <= _zz_12355[15 : 0];
        data_mid_119_imag <= _zz_12359[15 : 0];
        data_mid_55_real <= _zz_12363[15 : 0];
        data_mid_55_imag <= _zz_12367[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_120_real <= _zz_12377[15 : 0];
        data_mid_120_imag <= _zz_12381[15 : 0];
        data_mid_56_real <= _zz_12385[15 : 0];
        data_mid_56_imag <= _zz_12389[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_121_real <= _zz_12399[15 : 0];
        data_mid_121_imag <= _zz_12403[15 : 0];
        data_mid_57_real <= _zz_12407[15 : 0];
        data_mid_57_imag <= _zz_12411[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_122_real <= _zz_12421[15 : 0];
        data_mid_122_imag <= _zz_12425[15 : 0];
        data_mid_58_real <= _zz_12429[15 : 0];
        data_mid_58_imag <= _zz_12433[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_123_real <= _zz_12443[15 : 0];
        data_mid_123_imag <= _zz_12447[15 : 0];
        data_mid_59_real <= _zz_12451[15 : 0];
        data_mid_59_imag <= _zz_12455[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_124_real <= _zz_12465[15 : 0];
        data_mid_124_imag <= _zz_12469[15 : 0];
        data_mid_60_real <= _zz_12473[15 : 0];
        data_mid_60_imag <= _zz_12477[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_125_real <= _zz_12487[15 : 0];
        data_mid_125_imag <= _zz_12491[15 : 0];
        data_mid_61_real <= _zz_12495[15 : 0];
        data_mid_61_imag <= _zz_12499[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_126_real <= _zz_12509[15 : 0];
        data_mid_126_imag <= _zz_12513[15 : 0];
        data_mid_62_real <= _zz_12517[15 : 0];
        data_mid_62_imag <= _zz_12521[15 : 0];
      end
      if((current_level_cnt_value == 3'b111))begin
        data_mid_127_real <= _zz_12531[15 : 0];
        data_mid_127_imag <= _zz_12535[15 : 0];
        data_mid_63_real <= _zz_12539[15 : 0];
        data_mid_63_imag <= _zz_12543[15 : 0];
      end
    end
    current_level_cnt_willOverflow_regNext <= current_level_cnt_willOverflow;
  end

  always @ (posedge clk or posedge reset) begin
    if (reset) begin
      current_level_cnt_value <= 3'b000;
      current_level_cond_period_minus_1 <= 1'b0;
    end else begin
      current_level_cnt_value <= current_level_cnt_valueNext;
      if(io_data_in_valid_regNext)begin
        current_level_cond_period_minus_1 <= 1'b1;
      end else begin
        if(current_level_cnt_willOverflow)begin
          current_level_cond_period_minus_1 <= 1'b0;
        end
      end
    end
  end


endmodule

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

module SInt32fixTo23_8_ROUNDTOINF (
  input      [31:0]   din,
  output     [15:0]   dout
);
  wire       [32:0]   _zz_9;
  wire       [32:0]   _zz_10;
  wire       [7:0]    _zz_11;
  wire       [24:0]   _zz_12;
  wire       [24:0]   _zz_13;
  wire       [32:0]   _zz_14;
  wire       [32:0]   _zz_15;
  wire       [32:0]   _zz_16;
  wire       [9:0]    _zz_17;
  wire       [8:0]    _zz_18;
  reg        [24:0]   _zz_1;
  wire       [31:0]   _zz_2;
  wire       [31:0]   _zz_3;
  wire       [31:0]   _zz_4;
  wire       [32:0]   _zz_5;
  wire       [31:0]   _zz_6;
  reg        [24:0]   _zz_7;
  reg        [15:0]   _zz_8;

  assign _zz_9 = {_zz_4[31],_zz_4};
  assign _zz_10 = {_zz_3[31],_zz_3};
  assign _zz_11 = _zz_5[7 : 0];
  assign _zz_12 = _zz_5[32 : 8];
  assign _zz_13 = 25'h0000001;
  assign _zz_14 = ($signed(_zz_15) + $signed(_zz_16));
  assign _zz_15 = {_zz_6[31],_zz_6};
  assign _zz_16 = {_zz_2[31],_zz_2};
  assign _zz_17 = _zz_1[24 : 15];
  assign _zz_18 = _zz_1[23 : 15];
  assign _zz_2 = {{24'h0,1'b1},7'h0};
  assign _zz_3 = {25'h1ffffff,7'h0};
  assign _zz_4 = din[31 : 0];
  assign _zz_5 = ($signed(_zz_9) + $signed(_zz_10));
  assign _zz_6 = din[31 : 0];
  always @ (*) begin
    if((_zz_11 != 8'h0))begin
      _zz_7 = ($signed(_zz_12) + $signed(_zz_13));
    end else begin
      _zz_7 = _zz_5[32 : 8];
    end
  end

  always @ (*) begin
    if(_zz_5[32])begin
      _zz_1 = _zz_7;
    end else begin
      _zz_1 = (_zz_14 >>> 8);
    end
  end

  always @ (*) begin
    if(_zz_1[24])begin
      if((! (_zz_17 == 10'h3ff)))begin
        _zz_8 = 16'h8000;
      end else begin
        _zz_8 = _zz_1[15 : 0];
      end
    end else begin
      if((_zz_18 != 9'h0))begin
        _zz_8 = 16'h7fff;
      end else begin
        _zz_8 = _zz_1[15 : 0];
      end
    end
  end

  assign dout = _zz_8;

endmodule
